MACRO INVx8_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX8_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.10700000 0.27900000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.31500000 0.06300000 0.44100000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.44100000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx8_ASAP7_75t_L
MACRO XNOR2xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XNOR2XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
        RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.36000000 0.20700000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.28800000 0.12500000 0.30600000 0.14400000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
        RECT 0.45000000 0.04500000 0.46800000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.46800000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.01800000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.11700000 0.24300000 ;
  END

END XNOR2xp5_ASAP7_75t_L
MACRO AO221x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO221X1_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B2

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.47700000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
        RECT 0.47700000 0.18900000 0.52200000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.42300000 0.08100000 0.44100000 0.10700000 ;
      RECT 0.42300000 0.10700000 0.46800000 0.12500000 ;
      RECT 0.45000000 0.12500000 0.46800000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.11700000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.17100000 0.24300000 ;
      RECT 0.20700000 0.22500000 0.33300000 0.24300000 ;
  END

END AO221x1_ASAP7_75t_L
MACRO AND2x6_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND2X6_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.25200000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.14400000 ;
        RECT 0.23400000 0.04500000 0.25200000 0.14400000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.54900000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.34200000 0.18900000 0.54900000 0.20700000 ;
        RECT 0.34200000 0.20700000 0.36000000 0.22500000 ;
        RECT 0.31500000 0.22500000 0.36000000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.30600000 0.20700000 ;
  END

END AND2x6_ASAP7_75t_L
MACRO A2O1A1Ixp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN A2O1A1IXP33_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.04500000 0.18900000 0.17100000 0.20700000 ;
  END

END A2O1A1Ixp33_ASAP7_75t_L
MACRO AOI221xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI221XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B2

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END A2

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.17100000 0.24300000 ;
  END

END AOI221xp5_ASAP7_75t_L
MACRO NOR2xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR2XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.216 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.21600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.21600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.02700000 0.19800000 0.04500000 ;
        RECT 0.18000000 0.04500000 0.19800000 0.18900000 ;
        RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B

  OBS

  END

END NOR2xp33_ASAP7_75t_L
MACRO OR4x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR4X1_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.02700000 0.06300000 0.04500000 ;
        RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
    END
  END Y

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.07200000 0.06300000 0.36000000 0.08100000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
      RECT 0.31500000 0.18900000 0.36000000 0.20700000 ;
  END

END OR4x1_ASAP7_75t_L
MACRO AND5x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND5X2_ASAP7_75T_L 0 0 ;
 SIZE  1.08 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.08000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.08000000 0.27900000 ;
    END
  END VDD

  PIN E
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END E

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.12600000 0.63000000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.72000000 0.12600000 0.73800000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.96300000 0.06300000 1.00800000 0.08100000 ;
        RECT 0.99000000 0.08100000 1.00800000 0.18900000 ;
        RECT 0.96300000 0.18900000 1.00800000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.58500000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.42300000 0.06300000 0.65700000 0.08100000 ;
      RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.10700000 ;
      RECT 0.77400000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.93600000 0.12500000 0.95400000 0.14400000 ;
      RECT 0.77400000 0.12500000 0.79200000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.79200000 0.20700000 ;
  END

END AND5x2_ASAP7_75t_L
MACRO OAI21xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI21XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.17100000 0.20700000 ;
    END
  END Y

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.17100000 0.04500000 ;
  END

END OAI21xp5_ASAP7_75t_L
MACRO OA333x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA333X1_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
        RECT 0.01800000 0.22500000 0.06300000 0.24300000 ;
    END
  END Y

  PIN C3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END C3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END B3

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.31500000 0.02700000 0.54900000 0.04500000 ;
      RECT 0.15300000 0.06300000 0.38700000 0.08100000 ;
      RECT 0.47700000 0.06300000 0.63000000 0.08100000 ;
      RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
      RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
      RECT 0.07200000 0.18900000 0.63000000 0.20700000 ;
  END

END OA333x1_ASAP7_75t_L
MACRO OA333x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA333X2_ASAP7_75T_L 0 0 ;
 SIZE  0.7020000000000001 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.70200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.70200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.07200000 0.22500000 0.11700000 0.24300000 ;
    END
  END Y

  PIN C3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END C1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END B3

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.10700000 0.52200000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.12600000 0.63000000 0.16300000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.36900000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.20700000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.53100000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.68400000 0.20700000 ;
  END

END OA333x2_ASAP7_75t_L
MACRO SDFHx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFHX3_ASAP7_75T_L 0 0 ;
 SIZE  1.4580000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.45800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.45800000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END D

  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END SI

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.84600000 0.06300000 0.98100000 0.08100000 ;
        RECT 0.28800000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
       LAYER M2 ;
        RECT 0.31300000 0.06300000 0.86600000 0.08100000 ;
       LAYER V1 ;
        RECT 0.31300000 0.06300000 0.33100000 0.08100000 ;
        RECT 0.84800000 0.06300000 0.86600000 0.08100000 ;
    END
  END SE

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.28700000 0.06300000 1.41300000 0.08100000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.22500000 ;
        RECT 1.28700000 0.22500000 1.41300000 0.24300000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.49500000 0.08100000 ;
      RECT 0.82800000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.55800000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.10700000 ;
      RECT 0.50200000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 1.19700000 0.06300000 1.23700000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.14500000 ;
      RECT 0.33200000 0.14500000 0.37000000 0.16300000 ;
      RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.10700000 ;
      RECT 0.18000000 0.10700000 0.25200000 0.12500000 ;
      RECT 0.18000000 0.12500000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.26100000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.82800000 0.14500000 0.90000000 0.16300000 ;
      RECT 0.82800000 0.16300000 0.84600000 0.18900000 ;
      RECT 0.81900000 0.18900000 0.85900000 0.20700000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.18900000 ;
      RECT 1.20400000 0.18900000 1.27800000 0.20700000 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.09000000 0.20700000 ;
      RECT 0.07200000 0.20700000 0.09000000 0.22500000 ;
      RECT 0.07200000 0.22500000 0.27900000 0.24300000 ;
      RECT 0.31500000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.68400000 0.20700000 ;
      RECT 0.53100000 0.20700000 0.54900000 0.22500000 ;
      RECT 0.47500000 0.22500000 0.54900000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.73800000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.22500000 ;
      RECT 0.77400000 0.22500000 0.86400000 0.24300000 ;
      RECT 0.85500000 0.02700000 1.03500000 0.04500000 ;
      RECT 1.01700000 0.04500000 1.03500000 0.10700000 ;
      RECT 0.99000000 0.10700000 1.06200000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.18900000 ;
      RECT 0.93600000 0.18900000 1.06200000 0.20700000 ;
      RECT 0.93600000 0.20700000 0.95400000 0.22500000 ;
      RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
      RECT 1.07100000 0.02700000 1.11600000 0.04500000 ;
      RECT 1.09800000 0.04500000 1.11600000 0.14500000 ;
      RECT 1.04400000 0.14500000 1.11600000 0.16300000 ;
      RECT 1.09800000 0.16300000 1.11600000 0.22500000 ;
      RECT 1.07100000 0.22500000 1.11600000 0.24300000 ;
      RECT 1.15200000 0.02700000 1.23100000 0.04500000 ;
      RECT 1.15200000 0.04500000 1.17000000 0.22500000 ;
      RECT 1.15200000 0.22500000 1.22600000 0.24300000 ;
     LAYER M2 ;
      RECT 0.96100000 0.06300000 1.22400000 0.08100000 ;
      RECT 0.23200000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 1.17000000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.84600000 0.20700000 ;
      RECT 1.04200000 0.18900000 1.22400000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.49500000 0.24300000 ;
     LAYER V1 ;
      RECT 0.96100000 0.06300000 0.97900000 0.08100000 ;
      RECT 1.20600000 0.06300000 1.22400000 0.08100000 ;
      RECT 0.23200000 0.10700000 0.25000000 0.12500000 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.84800000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 0.36000000 0.16300000 ;
      RECT 1.15200000 0.14500000 1.17000000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.68200000 0.20700000 ;
      RECT 0.82800000 0.18900000 0.84600000 0.20700000 ;
      RECT 1.04200000 0.18900000 1.06000000 0.20700000 ;
      RECT 1.20600000 0.18900000 1.22400000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.27700000 0.24300000 ;
      RECT 0.47700000 0.22500000 0.49500000 0.24300000 ;
  END

END SDFHx3_ASAP7_75t_L
MACRO INVx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX2_ASAP7_75T_L 0 0 ;
 SIZE  0.216 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.21600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.21600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx2_ASAP7_75t_L
MACRO AO332x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO332X2_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.12600000 0.06300000 0.63000000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.63000000 0.20700000 ;
      RECT 0.36900000 0.22500000 0.60300000 0.24300000 ;
  END

END AO332x2_ASAP7_75t_L
MACRO OAI32xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI32XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.04500000 0.18900000 0.36000000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
  END

END OAI32xp33_ASAP7_75t_L
MACRO CKINVDCx6p67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX6P67_ASAP7_75T_L 0 0 ;
 SIZE  1.296 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.29600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.29600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.34000000 0.10700000 0.52200000 0.12500000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
       LAYER M2 ;
        RECT 0.17800000 0.10700000 0.36000000 0.12500000 ;
       LAYER V1 ;
        RECT 0.17800000 0.10700000 0.19600000 0.12500000 ;
        RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.76500000 0.04500000 ;
        RECT 1.07100000 0.06300000 1.19700000 0.08100000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.14400000 0.20700000 ;
        RECT 0.12600000 0.20700000 0.14400000 0.22500000 ;
        RECT 1.09800000 0.08100000 1.11600000 0.22500000 ;
        RECT 0.12600000 0.22500000 1.19700000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.53100000 0.06300000 0.65700000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.14400000 ;
      RECT 0.85500000 0.06300000 0.98100000 0.08100000 ;
      RECT 0.93600000 0.08100000 0.95400000 0.14400000 ;
      RECT 0.80100000 0.02700000 1.03500000 0.04500000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.10700000 ;
      RECT 1.01700000 0.04500000 1.03500000 0.10700000 ;
      RECT 0.66400000 0.10700000 0.81900000 0.12500000 ;
      RECT 1.01700000 0.10700000 1.06200000 0.12500000 ;
      RECT 0.72000000 0.12500000 0.73800000 0.14400000 ;
      RECT 1.04400000 0.12500000 1.06200000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.85500000 0.18900000 0.98100000 0.20700000 ;
     LAYER M2 ;
      RECT 0.50200000 0.10700000 0.68400000 0.12500000 ;
     LAYER V1 ;
      RECT 0.50200000 0.10700000 0.52000000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
  END

END CKINVDCx6p67_ASAP7_75t_L
MACRO AOI211xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI211XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.22500000 0.17100000 0.24300000 ;
  END

END AOI211xp5_ASAP7_75t_L
MACRO MAJx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN MAJX2_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.27900000 0.08100000 ;
        RECT 0.15300000 0.08100000 0.17100000 0.10700000 ;
        RECT 0.26100000 0.08100000 0.27900000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.17100000 0.12500000 ;
        RECT 0.26100000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.28800000 0.12500000 0.30600000 0.14400000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.12600000 0.22500000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.36900000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.22500000 ;
        RECT 0.36900000 0.22500000 0.41400000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END MAJx2_ASAP7_75t_L
MACRO AOI322xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI322XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.36900000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.18900000 0.27900000 0.20700000 ;
      RECT 0.20700000 0.22500000 0.44100000 0.24300000 ;
  END

END AOI322xp5_ASAP7_75t_L
MACRO AND2x4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND2X4_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.22500000 0.04500000 ;
        RECT 0.20700000 0.04500000 0.22500000 0.06300000 ;
        RECT 0.20700000 0.06300000 0.25200000 0.08100000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.14400000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.44100000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.34200000 0.18900000 0.44100000 0.20700000 ;
        RECT 0.34200000 0.20700000 0.36000000 0.22500000 ;
        RECT 0.31500000 0.22500000 0.36000000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.12600000 0.06300000 0.17100000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.30600000 0.20700000 ;
  END

END AND2x4_ASAP7_75t_L
MACRO TIEHIx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN TIEHIX1_ASAP7_75T_L 0 0 ;
 SIZE  0.16200000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.16200000 0.27900000 ;
    END
  END VDD

  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.16200000 0.00900000 ;
    END
  END VSS

  PIN H
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.06700000 0.07000000 0.14400000 0.08800000 ;
        RECT 0.12600000 0.08800000 0.14400000 0.22500000 ;
        RECT 0.09400000 0.22500000 0.14400000 0.24300000 ;
    END
  END H

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.02700000 0.06800000 0.04500000 ;
      RECT 0.01800000 0.04500000 0.03600000 0.15500000 ;
      RECT 0.01800000 0.15500000 0.09500000 0.17300000 ;
  END

END TIEHIx1_ASAP7_75t_L
MACRO DECAPx6_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DECAPX6_ASAP7_75T_L 0 0 ;
 SIZE  0.756 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.75600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.75600000 0.27900000 ;
    END
  END VDD

  OBS
     LAYER M1 ;
      RECT 0.34200000 0.06300000 0.71100000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.41400000 0.20700000 ;
  END

END DECAPx6_ASAP7_75t_L
MACRO OA331x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA331X2_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.07200000 0.22500000 0.11700000 0.24300000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.14400000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B3

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.10700000 0.52200000 0.14400000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.36900000 0.06300000 0.49500000 0.08100000 ;
      RECT 0.53100000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.57600000 0.20700000 ;
  END

END OA331x2_ASAP7_75t_L
MACRO BUFx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX4_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.27900000 0.04500000 ;
        RECT 0.26100000 0.04500000 0.27900000 0.22500000 ;
        RECT 0.15300000 0.22500000 0.27900000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx4_ASAP7_75t_L
MACRO HB2xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HB2XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.25200000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.25200000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.09000000 0.04500000 ;
      RECT 0.07200000 0.04500000 0.09000000 0.06300000 ;
      RECT 0.07200000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14500000 ;
      RECT 0.18000000 0.12600000 0.19800000 0.14500000 ;
      RECT 0.12600000 0.14500000 0.19800000 0.16300000 ;
      RECT 0.12600000 0.16300000 0.14400000 0.22500000 ;
      RECT 0.04500000 0.22500000 0.14400000 0.24300000 ;
  END

END HB2xp67_ASAP7_75t_L
MACRO BUFx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX2_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
        RECT 0.18000000 0.04500000 0.19800000 0.18900000 ;
        RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
  END

END BUFx2_ASAP7_75t_L
MACRO DHLx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DHLX2_ASAP7_75T_L 0 0 ;
 SIZE  0.8640000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.86400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.86400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
        RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
        RECT 0.74700000 0.18900000 0.79200000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.66400000 0.10700000 0.73800000 0.12500000 ;
      RECT 0.72000000 0.12500000 0.73800000 0.14400000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.16400000 ;
      RECT 0.09900000 0.02700000 0.36000000 0.04500000 ;
      RECT 0.09900000 0.04500000 0.11700000 0.06300000 ;
      RECT 0.34200000 0.04500000 0.36000000 0.06300000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.34200000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.41400000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.42300000 0.02700000 0.54900000 0.04500000 ;
      RECT 0.53100000 0.04500000 0.54900000 0.06300000 ;
      RECT 0.53100000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.50400000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.50400000 0.20700000 0.52200000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.58500000 0.02700000 0.63000000 0.04500000 ;
      RECT 0.61200000 0.04500000 0.63000000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.63000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.55800000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.63000000 0.16200000 ;
     LAYER V1 ;
      RECT 0.55800000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.52200000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
  END

END DHLx2_ASAP7_75t_L
MACRO DLLx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DLLX1_ASAP7_75T_L 0 0 ;
 SIZE  0.8100000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.81000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.81000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
        RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
        RECT 0.74700000 0.18900000 0.79200000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.66400000 0.10700000 0.73800000 0.12500000 ;
      RECT 0.72000000 0.12500000 0.73800000 0.14400000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.16400000 ;
      RECT 0.01800000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.06300000 ;
      RECT 0.45000000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.50400000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.50400000 0.20700000 0.52200000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.58500000 0.02700000 0.63000000 0.04500000 ;
      RECT 0.61200000 0.04500000 0.63000000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.63000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.55800000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.63000000 0.16200000 ;
     LAYER V1 ;
      RECT 0.55800000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.52200000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
  END

END DLLx1_ASAP7_75t_L
MACRO NOR2x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR2X2_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.14500000 ;
        RECT 0.39600000 0.12600000 0.41400000 0.14500000 ;
        RECT 0.12600000 0.14500000 0.17100000 0.16300000 ;
        RECT 0.36900000 0.14500000 0.41400000 0.16300000 ;
        RECT 0.15300000 0.16300000 0.17100000 0.18900000 ;
        RECT 0.36900000 0.16300000 0.38700000 0.18900000 ;
        RECT 0.15300000 0.18900000 0.38700000 0.20700000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
        RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.12600000 0.27900000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.22500000 0.49500000 0.24300000 ;
  END

END NOR2x2_ASAP7_75t_L
MACRO DECAPx2b_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DECAPX2B_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.18000000 0.12600000 0.19800000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
  END

END DECAPx2b_ASAP7_75t_L
MACRO DFFHQNx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFHQNX3_ASAP7_75T_L 0 0 ;
 SIZE  1.1880000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.18800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.18800000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.01700000 0.06300000 1.14300000 0.08100000 ;
        RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
        RECT 1.01700000 0.18900000 1.14300000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.08300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.08300000 ;
      RECT 0.66600000 0.10500000 0.68400000 0.14400000 ;
      RECT 0.93600000 0.06100000 0.95400000 0.10700000 ;
      RECT 0.93600000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.16400000 ;
      RECT 0.01800000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.54800000 0.06300000 0.58600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.55000000 0.18900000 0.58700000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.39600000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.39600000 0.20700000 0.41400000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.41400000 0.24300000 ;
      RECT 0.50400000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.50400000 0.22500000 0.54100000 0.24300000 ;
      RECT 0.58000000 0.22500000 0.62800000 0.24300000 ;
      RECT 0.81800000 0.06300000 0.85500000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.90000000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.45000000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.72000000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.58600000 0.20700000 ;
      RECT 0.51200000 0.22500000 0.62700000 0.24300000 ;
     LAYER V1 ;
      RECT 0.45000000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.55800000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.72000000 0.06300000 0.73800000 0.08100000 ;
      RECT 0.82800000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.93600000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.36000000 0.16200000 ;
      RECT 0.45000000 0.14400000 0.46800000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.46600000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.52100000 0.22500000 0.53900000 0.24300000 ;
      RECT 0.59300000 0.22500000 0.61100000 0.24300000 ;
  END

END DFFHQNx3_ASAP7_75t_L
MACRO AOI31xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI31XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.7020000000000001 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.70200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.70200000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A3

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.25200000 0.08100000 ;
        RECT 0.47700000 0.06300000 0.54900000 0.08100000 ;
        RECT 0.47700000 0.08100000 0.49500000 0.10700000 ;
        RECT 0.45000000 0.10700000 0.49500000 0.12500000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.45000000 0.12500000 0.46800000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.36900000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
      RECT 0.31500000 0.04500000 0.33300000 0.06300000 ;
      RECT 0.31500000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.04500000 0.22500000 0.54900000 0.24300000 ;
  END

END AOI31xp67_ASAP7_75t_L
MACRO OA332x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA332X1_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
        RECT 0.01800000 0.22500000 0.06300000 0.24300000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END B3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.31500000 0.02700000 0.54900000 0.04500000 ;
      RECT 0.15300000 0.06300000 0.38700000 0.08100000 ;
      RECT 0.47700000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.07200000 0.18900000 0.57600000 0.20700000 ;
  END

END OA332x1_ASAP7_75t_L
MACRO AND3x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND3X1_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.30600000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.23400000 0.12600000 0.25200000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.25200000 0.20700000 ;
  END

END AND3x1_ASAP7_75t_L
MACRO CKINVDCx10_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX10_ASAP7_75T_L 0 0 ;
 SIZE  1.296 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.29600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.29600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.34000000 0.10700000 0.52200000 0.12500000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
       LAYER M2 ;
        RECT 0.17800000 0.10700000 0.36000000 0.12500000 ;
       LAYER V1 ;
        RECT 0.17800000 0.10700000 0.19600000 0.12500000 ;
        RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.76500000 0.04500000 ;
        RECT 1.07100000 0.06300000 1.19700000 0.08100000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.14400000 0.20700000 ;
        RECT 0.12600000 0.20700000 0.14400000 0.22500000 ;
        RECT 1.09800000 0.08100000 1.11600000 0.22500000 ;
        RECT 0.12600000 0.22500000 1.19700000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.53100000 0.06300000 0.65700000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.14400000 ;
      RECT 0.85500000 0.06300000 0.98100000 0.08100000 ;
      RECT 0.93600000 0.08100000 0.95400000 0.14400000 ;
      RECT 0.80100000 0.02700000 1.03500000 0.04500000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.10700000 ;
      RECT 1.01700000 0.04500000 1.03500000 0.10700000 ;
      RECT 0.66400000 0.10700000 0.81900000 0.12500000 ;
      RECT 1.01700000 0.10700000 1.06200000 0.12500000 ;
      RECT 0.72000000 0.12500000 0.73800000 0.14400000 ;
      RECT 1.04400000 0.12500000 1.06200000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.85500000 0.18900000 0.98100000 0.20700000 ;
     LAYER M2 ;
      RECT 0.50200000 0.10700000 0.68400000 0.12500000 ;
     LAYER V1 ;
      RECT 0.50200000 0.10700000 0.52000000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
  END

END CKINVDCx10_ASAP7_75t_L
MACRO ICGx5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX5_ASAP7_75T_L 0 0 ;
 SIZE  1.1880000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.18800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.18800000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END SE

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.06300000 0.73800000 0.08100000 ;
        RECT 0.72000000 0.08100000 0.73800000 0.14400000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.16500000 ;
        RECT 0.23400000 0.12600000 0.25200000 0.18900000 ;
        RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
        RECT 0.23400000 0.18900000 0.36000000 0.20700000 ;
       LAYER M2 ;
        RECT 0.34200000 0.14500000 0.63000000 0.16300000 ;
       LAYER V1 ;
        RECT 0.34200000 0.14500000 0.36000000 0.16300000 ;
        RECT 0.61200000 0.14500000 0.63000000 0.16300000 ;
    END
  END CLK

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.90900000 0.02700000 0.95400000 0.04500000 ;
        RECT 0.93600000 0.04500000 0.95400000 0.06300000 ;
        RECT 0.93600000 0.06300000 1.14300000 0.08100000 ;
        RECT 0.93600000 0.08100000 0.95400000 0.18900000 ;
        RECT 0.93600000 0.18900000 1.14300000 0.20700000 ;
        RECT 0.93600000 0.20700000 0.95400000 0.22500000 ;
        RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
    END
  END GCLK

  OBS
     LAYER M1 ;
      RECT 0.28800000 0.06300000 0.38700000 0.08100000 ;
      RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
      RECT 0.39600000 0.10500000 0.41400000 0.14400000 ;
      RECT 0.09900000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.55800000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.55800000 0.04500000 0.57600000 0.18900000 ;
      RECT 0.55800000 0.18900000 0.60300000 0.20700000 ;
      RECT 0.31500000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.42300000 0.04500000 0.44100000 0.06300000 ;
      RECT 0.42300000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
      RECT 0.38600000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.38600000 0.20700000 0.40400000 0.22500000 ;
      RECT 0.26100000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.47700000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.47700000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.82800000 0.12600000 0.84600000 0.14500000 ;
      RECT 0.80100000 0.14500000 0.84600000 0.16300000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.18900000 ;
      RECT 0.80100000 0.16300000 0.81900000 0.18900000 ;
      RECT 0.63900000 0.18900000 0.81900000 0.20700000 ;
      RECT 0.63900000 0.20700000 0.65700000 0.22500000 ;
      RECT 0.55600000 0.22500000 0.65700000 0.24300000 ;
      RECT 0.74700000 0.02700000 0.79200000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.06300000 ;
      RECT 0.77400000 0.06300000 0.90000000 0.08100000 ;
      RECT 0.88200000 0.08100000 0.90000000 0.18900000 ;
      RECT 0.85500000 0.18900000 0.90000000 0.20700000 ;
      RECT 0.85500000 0.20700000 0.87300000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.87300000 0.24300000 ;
     LAYER M2 ;
      RECT 0.36000000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.42100000 0.22500000 0.57600000 0.24300000 ;
     LAYER V1 ;
      RECT 0.36600000 0.06300000 0.38400000 0.08100000 ;
      RECT 0.55800000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.42100000 0.22500000 0.43900000 0.24300000 ;
      RECT 0.55800000 0.22500000 0.57600000 0.24300000 ;
  END

END ICGx5_ASAP7_75t_L
MACRO OA332x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA332X2_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.07200000 0.22500000 0.11700000 0.24300000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END B3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.10700000 0.52200000 0.14400000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.36900000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.20700000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.53100000 0.06300000 0.63000000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.63000000 0.20700000 ;
  END

END OA332x2_ASAP7_75t_L
MACRO DECAPx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DECAPX1_ASAP7_75T_L 0 0 ;
 SIZE  0.216 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.21600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.21600000 0.27900000 ;
    END
  END VDD

  OBS
     LAYER M1 ;
      RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
  END

END DECAPx1_ASAP7_75t_L
MACRO FAx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN FAX1_ASAP7_75T_L 0 0 ;
 SIZE  0.7560000000000006 BY 0.2700000000000002 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN SN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.35500000 0.02700000 0.49500000 0.04500000 ;
        RECT 0.35500000 0.04500000 0.37400000 0.18900000 ;
        RECT 0.35500000 0.18900000 0.49500000 0.20700000 ;
    END
  END SN

  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.75600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.75600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10500000 0.09000000 0.14400000 ;
        RECT 0.61200000 0.10500000 0.63000000 0.14400000 ;
        RECT 0.39600000 0.10500000 0.41400000 0.16300000 ;
       LAYER M2 ;
        RECT 0.07200000 0.10700000 0.63000000 0.12500000 ;
       LAYER V1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.12500000 ;
        RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.66600000 0.12600000 0.68400000 0.14500000 ;
        RECT 0.66600000 0.14500000 0.71100000 0.16300000 ;
        RECT 0.18000000 0.12600000 0.19800000 0.18800000 ;
        RECT 0.31900000 0.12600000 0.33700000 0.18800000 ;
        RECT 0.18000000 0.18800000 0.33700000 0.20600000 ;
        RECT 0.31900000 0.20600000 0.33700000 0.22500000 ;
        RECT 0.69300000 0.16300000 0.71100000 0.22500000 ;
        RECT 0.31900000 0.22500000 0.71100000 0.24300000 ;
    END
  END B

  PIN CON
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42100000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.14400000 ;
        RECT 0.12600000 0.06300000 0.33000000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.22500000 ;
        RECT 0.12600000 0.22500000 0.22400000 0.24300000 ;
       LAYER M2 ;
        RECT 0.31000000 0.06300000 0.44100000 0.08100000 ;
       LAYER V1 ;
        RECT 0.31000000 0.06300000 0.32800000 0.08100000 ;
        RECT 0.42300000 0.06300000 0.44100000 0.08100000 ;
    END
  END CON

  PIN CI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.14500000 ;
        RECT 0.23400000 0.14500000 0.27900000 0.16300000 ;
        RECT 0.45000000 0.12600000 0.46800000 0.14500000 ;
        RECT 0.44100000 0.14500000 0.47700000 0.16300000 ;
        RECT 0.55800000 0.12600000 0.57600000 0.14500000 ;
        RECT 0.54900000 0.14500000 0.58500000 0.16300000 ;
       LAYER M2 ;
        RECT 0.25900000 0.14500000 0.57600000 0.16300000 ;
       LAYER V1 ;
        RECT 0.25900000 0.14500000 0.27700000 0.16300000 ;
        RECT 0.45000000 0.14500000 0.46800000 0.16300000 ;
        RECT 0.55800000 0.14500000 0.57600000 0.16300000 ;
    END
  END CI

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.53100000 0.02700000 0.65700000 0.04500000 ;
      RECT 0.53100000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.09000000 0.24300000 ;
      RECT 0.25600000 0.22500000 0.29300000 0.24300000 ;
     LAYER M2 ;
      RECT 0.07000000 0.22500000 0.27900000 0.24300000 ;
     LAYER V1 ;
      RECT 0.07000000 0.22500000 0.08800000 0.24300000 ;
      RECT 0.26100000 0.22500000 0.27900000 0.24300000 ;
  END

END FAx1_ASAP7_75t_L
MACRO AOI311xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI311XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.31500000 0.18900000 0.36000000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
  END

END AOI311xp33_ASAP7_75t_L
MACRO OAI321xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI321XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END C

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
  END

END OAI321xp33_ASAP7_75t_L
MACRO OR3x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR3X2_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.30600000 0.04500000 ;
        RECT 0.28800000 0.04500000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
  END

END OR3x2_ASAP7_75t_L
MACRO BUFx16f_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX16F_ASAP7_75T_L 0 0 ;
 SIZE  1.188 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.18800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.18800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 1.08900000 0.08100000 ;
        RECT 0.36900000 0.08100000 0.38700000 0.18900000 ;
        RECT 0.31500000 0.18900000 1.08900000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.10700000 ;
      RECT 0.23400000 0.10700000 0.30600000 0.12500000 ;
      RECT 0.28800000 0.12500000 0.30600000 0.14400000 ;
      RECT 0.23400000 0.12500000 0.25200000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.25200000 0.20700000 ;
  END

END BUFx16f_ASAP7_75t_L
MACRO AND3x4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND3X4_ASAP7_75T_L 0 0 ;
 SIZE  0.756 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.75600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.75600000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.53100000 0.12600000 0.54900000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.66600000 0.12600000 0.68400000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.47700000 0.02700000 0.71100000 0.04500000 ;
      RECT 0.31500000 0.06300000 0.54900000 0.08100000 ;
      RECT 0.61200000 0.06300000 0.65700000 0.08100000 ;
      RECT 0.23400000 0.12600000 0.25200000 0.14500000 ;
      RECT 0.23400000 0.14500000 0.27900000 0.16300000 ;
      RECT 0.26100000 0.16300000 0.27900000 0.18900000 ;
      RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
      RECT 0.26100000 0.18900000 0.65700000 0.20700000 ;
  END

END AND3x4_ASAP7_75t_L
MACRO OAI33xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI33XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A3

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
  END

END OAI33xp33_ASAP7_75t_L
MACRO INVx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX1_ASAP7_75T_L 0 0 ;
 SIZE  0.162 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.16200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.16200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  OBS

  END

END INVx1_ASAP7_75t_L
MACRO DLLx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DLLX2_ASAP7_75T_L 0 0 ;
 SIZE  0.8640000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.86400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.86400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.69300000 0.06300000 0.81900000 0.08100000 ;
        RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
        RECT 0.69300000 0.18900000 0.81900000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.66400000 0.10700000 0.73800000 0.12500000 ;
      RECT 0.72000000 0.12500000 0.73800000 0.14400000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.16400000 ;
      RECT 0.07200000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.07200000 0.04500000 0.09000000 0.06300000 ;
      RECT 0.26100000 0.04500000 0.27900000 0.06300000 ;
      RECT 0.01800000 0.06300000 0.09000000 0.08100000 ;
      RECT 0.26100000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.42300000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.47700000 0.04500000 0.49500000 0.06300000 ;
      RECT 0.47700000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.50400000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.50400000 0.20700000 0.52200000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.58500000 0.02700000 0.63000000 0.04500000 ;
      RECT 0.61200000 0.04500000 0.63000000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.63000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.55800000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.63000000 0.16200000 ;
     LAYER V1 ;
      RECT 0.55800000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.52200000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
  END

END DLLx2_ASAP7_75t_L
MACRO MAJIxp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN MAJIXP5_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.14500000 ;
        RECT 0.23400000 0.12600000 0.25200000 0.14500000 ;
        RECT 0.07200000 0.14500000 0.11700000 0.16300000 ;
        RECT 0.20700000 0.14500000 0.25200000 0.16300000 ;
        RECT 0.09900000 0.16300000 0.11700000 0.18900000 ;
        RECT 0.20700000 0.16300000 0.22500000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.12600000 0.17100000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.36000000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
      RECT 0.09900000 0.22500000 0.33300000 0.24300000 ;
  END

END MAJIxp5_ASAP7_75t_L
MACRO HB1xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HB1XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.216 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.21600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.21600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
        RECT 0.18000000 0.04500000 0.19800000 0.22500000 ;
        RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.11700000 0.04500000 ;
      RECT 0.09900000 0.04500000 0.11700000 0.06300000 ;
      RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.09900000 0.20700000 0.11700000 0.22500000 ;
      RECT 0.04500000 0.22500000 0.11700000 0.24300000 ;
  END

END HB1xp67_ASAP7_75t_L
MACRO AO333x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO333X1_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.02700000 0.06300000 0.04500000 ;
        RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B3

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B1

  PIN C3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.07200000 0.06300000 0.63000000 0.08100000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
      RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
      RECT 0.47700000 0.18900000 0.63000000 0.20700000 ;
      RECT 0.31500000 0.22500000 0.54900000 0.24300000 ;
  END

END AO333x1_ASAP7_75t_L
MACRO XOR2x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XOR2X1_ASAP7_75T_L 0 0 ;
 SIZE  0.6480000000000001 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.14500000 ;
        RECT 0.47500000 0.14500000 0.52200000 0.16300000 ;
        RECT 0.34200000 0.12600000 0.36000000 0.14500000 ;
        RECT 0.34200000 0.14500000 0.38700000 0.16300000 ;
        RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
        RECT 0.34200000 0.16300000 0.36000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.36000000 0.20700000 ;
       LAYER M2 ;
        RECT 0.35800000 0.14500000 0.49500000 0.16300000 ;
       LAYER V1 ;
        RECT 0.36400000 0.14500000 0.38200000 0.16300000 ;
        RECT 0.47700000 0.14500000 0.49500000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.06300000 0.57600000 0.08100000 ;
        RECT 0.55800000 0.08100000 0.57600000 0.14400000 ;
        RECT 0.12600000 0.12600000 0.14400000 0.14500000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14500000 ;
        RECT 0.12600000 0.14500000 0.30600000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.63000000 0.04500000 ;
        RECT 0.61200000 0.04500000 0.63000000 0.18900000 ;
        RECT 0.42300000 0.18900000 0.63000000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.39400000 0.10700000 0.44100000 0.12500000 ;
      RECT 0.42300000 0.12500000 0.44100000 0.14400000 ;
      RECT 0.01800000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.10700000 ;
      RECT 0.18000000 0.10700000 0.25200000 0.12500000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.17100000 0.24300000 ;
      RECT 0.26100000 0.22500000 0.60300000 0.24300000 ;
     LAYER M2 ;
      RECT 0.23200000 0.10700000 0.42000000 0.12500000 ;
     LAYER V1 ;
      RECT 0.23200000 0.10700000 0.25000000 0.12500000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
  END

END XOR2x1_ASAP7_75t_L
MACRO OAI31xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI31XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.22500000 0.04500000 ;
  END

END OAI31xp33_ASAP7_75t_L
MACRO OAI31xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI31XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.7020000000000001 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.70200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.70200000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A3

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.14500000 ;
        RECT 0.45000000 0.14500000 0.52200000 0.16300000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.50400000 0.16300000 0.52200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.25200000 0.20700000 ;
        RECT 0.50400000 0.18900000 0.54900000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.10700000 0.57600000 0.14400000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.54900000 0.04500000 ;
      RECT 0.28800000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.28800000 0.20700000 0.30600000 0.22500000 ;
      RECT 0.09900000 0.22500000 0.30600000 0.24300000 ;
      RECT 0.36900000 0.22500000 0.60300000 0.24300000 ;
  END

END OAI31xp67_ASAP7_75t_L
MACRO OAI221xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI221XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B2

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END C

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END A2

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.17100000 0.04500000 ;
      RECT 0.20700000 0.02700000 0.33300000 0.04500000 ;
  END

END OAI221xp5_ASAP7_75t_L
MACRO OAI222xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI222XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.38700000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END C1

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END C2

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.20700000 0.06300000 0.44100000 0.08100000 ;
  END

END OAI222xp33_ASAP7_75t_L
MACRO CKINVDCx12_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX12_ASAP7_75T_L 0 0 ;
 SIZE  1.4040000000000001 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.40400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.40400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.38700000 0.04500000 ;
        RECT 0.15300000 0.04500000 0.17100000 0.10700000 ;
        RECT 0.36900000 0.04500000 0.38700000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.17100000 0.12500000 ;
        RECT 0.36900000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
        RECT 0.85500000 0.06300000 0.98100000 0.08100000 ;
        RECT 1.28700000 0.06300000 1.33200000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.22500000 ;
        RECT 0.88200000 0.08100000 0.90000000 0.22500000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.22500000 ;
        RECT 0.07200000 0.22500000 1.33200000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.63900000 0.06300000 0.76500000 0.08100000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 0.58500000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.58500000 0.04500000 0.60300000 0.10700000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.10700000 ;
      RECT 0.55800000 0.10700000 0.60300000 0.12500000 ;
      RECT 0.80100000 0.10700000 0.84600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.82800000 0.12500000 0.84600000 0.14400000 ;
      RECT 1.07100000 0.06300000 1.19700000 0.08100000 ;
      RECT 1.15200000 0.08100000 1.17000000 0.14400000 ;
      RECT 1.01700000 0.02700000 1.25100000 0.04500000 ;
      RECT 1.01700000 0.04500000 1.03500000 0.10700000 ;
      RECT 1.23300000 0.04500000 1.25100000 0.10700000 ;
      RECT 0.99000000 0.10700000 1.03500000 0.12500000 ;
      RECT 1.23300000 0.10700000 1.27800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 1.26000000 0.12500000 1.27800000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.63900000 0.18900000 0.76500000 0.20700000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.18900000 ;
      RECT 1.07100000 0.18900000 1.19700000 0.20700000 ;
  END

END CKINVDCx12_ASAP7_75t_L
MACRO DLLx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DLLX3_ASAP7_75T_L 0 0 ;
 SIZE  0.9180000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.91800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.91800000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.74700000 0.06300000 0.87300000 0.08100000 ;
        RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
        RECT 0.74700000 0.18900000 0.87300000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.50400000 0.10500000 0.52200000 0.14400000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.14500000 ;
      RECT 0.66400000 0.14500000 0.73800000 0.16300000 ;
      RECT 0.07200000 0.02700000 0.30600000 0.04500000 ;
      RECT 0.07200000 0.04500000 0.09000000 0.06300000 ;
      RECT 0.28800000 0.04500000 0.30600000 0.06300000 ;
      RECT 0.01800000 0.06300000 0.09000000 0.08100000 ;
      RECT 0.28800000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.42300000 0.02700000 0.54900000 0.04500000 ;
      RECT 0.53100000 0.04500000 0.54900000 0.06300000 ;
      RECT 0.53100000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.50400000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.50400000 0.20700000 0.52200000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.58500000 0.02700000 0.63000000 0.04500000 ;
      RECT 0.61200000 0.04500000 0.63000000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.63000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.50400000 0.10700000 0.63000000 0.12500000 ;
      RECT 0.55800000 0.14500000 0.68400000 0.16300000 ;
     LAYER V1 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
      RECT 0.55800000 0.14500000 0.57600000 0.16300000 ;
      RECT 0.66600000 0.14500000 0.68400000 0.16300000 ;
  END

END DLLx3_ASAP7_75t_L
MACRO NAND3x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND3X2_ASAP7_75T_L 0 0 ;
 SIZE  1.08 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.08000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.08000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.04500000 0.06300000 0.17100000 0.08100000 ;
        RECT 0.90900000 0.06300000 1.03500000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.22500000 ;
        RECT 0.93600000 0.08100000 0.95400000 0.22500000 ;
        RECT 0.12600000 0.22500000 0.95400000 0.24300000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.14500000 ;
        RECT 0.88200000 0.12600000 0.90000000 0.14500000 ;
        RECT 0.18000000 0.14500000 0.30600000 0.16300000 ;
        RECT 0.85500000 0.14500000 0.90000000 0.16300000 ;
        RECT 0.28800000 0.16300000 0.30600000 0.18900000 ;
        RECT 0.85500000 0.16300000 0.87300000 0.18900000 ;
        RECT 0.28800000 0.18900000 0.87300000 0.20700000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.06300000 0.63000000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.10700000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.10700000 ;
        RECT 0.34200000 0.10700000 0.52200000 0.12500000 ;
        RECT 0.61200000 0.10700000 0.73800000 0.12500000 ;
        RECT 0.34200000 0.12500000 0.36000000 0.14400000 ;
        RECT 0.72000000 0.12500000 0.73800000 0.14400000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
      RECT 0.74700000 0.02700000 0.98100000 0.04500000 ;
      RECT 0.45000000 0.02700000 0.68400000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.06300000 ;
      RECT 0.66600000 0.04500000 0.68400000 0.06300000 ;
      RECT 0.26100000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.66600000 0.06300000 0.81900000 0.08100000 ;
  END

END NAND3x2_ASAP7_75t_L
MACRO AOI21x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI21X1_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.02700000 0.41400000 0.04500000 ;
        RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
        RECT 0.39600000 0.04500000 0.41400000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
        RECT 0.36900000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
    END
  END B

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.14500000 ;
        RECT 0.26100000 0.14500000 0.30600000 0.16300000 ;
        RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
        RECT 0.26100000 0.16300000 0.27900000 0.18900000 ;
        RECT 0.12600000 0.18900000 0.27900000 0.20700000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.12600000 0.22500000 0.16300000 ;
    END
  END A2

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.22500000 0.33300000 0.24300000 ;
  END

END AOI21x1_ASAP7_75t_L
MACRO NAND2xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND2XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.216 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.21600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.21600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.19800000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B

  OBS

  END

END NAND2xp5_ASAP7_75t_L
MACRO NAND3xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND3XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.17100000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END C

  OBS

  END

END NAND3xp33_ASAP7_75t_L
MACRO BUFx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX3_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.27900000 0.04500000 ;
        RECT 0.20700000 0.04500000 0.22500000 0.18900000 ;
        RECT 0.18000000 0.18900000 0.27900000 0.20700000 ;
        RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
        RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx3_ASAP7_75t_L
MACRO AO331x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO331X2_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B3

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.36900000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.12600000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.20700000 0.22500000 0.44100000 0.24300000 ;
  END

END AO331x2_ASAP7_75t_L
MACRO INVx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX3_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx3_ASAP7_75t_L
MACRO CKINVDCx8_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX8_ASAP7_75T_L 0 0 ;
 SIZE  1.188 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.18800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.18800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.14500000 ;
        RECT 0.39600000 0.12600000 0.41400000 0.14500000 ;
        RECT 0.72000000 0.12600000 0.73800000 0.14500000 ;
        RECT 1.04400000 0.12600000 1.06200000 0.14500000 ;
        RECT 0.12600000 0.14500000 0.17100000 0.16300000 ;
        RECT 0.36900000 0.14500000 0.41400000 0.16300000 ;
        RECT 0.69300000 0.14500000 0.73800000 0.16300000 ;
        RECT 1.01700000 0.14500000 1.06200000 0.16300000 ;
        RECT 0.15300000 0.16300000 0.17100000 0.22500000 ;
        RECT 0.36900000 0.16300000 0.38700000 0.22500000 ;
        RECT 0.69300000 0.16300000 0.71100000 0.22500000 ;
        RECT 1.01700000 0.16300000 1.03500000 0.22500000 ;
        RECT 0.15300000 0.22500000 1.03500000 0.24300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 1.06200000 0.04500000 ;
        RECT 0.15300000 0.04500000 0.17100000 0.06300000 ;
        RECT 1.04400000 0.04500000 1.06200000 0.06300000 ;
        RECT 0.07200000 0.06300000 0.17100000 0.08100000 ;
        RECT 1.04400000 0.06300000 1.11600000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.45000000 0.04500000 0.46800000 0.18900000 ;
        RECT 0.77400000 0.04500000 0.79200000 0.18900000 ;
        RECT 1.09800000 0.08100000 1.11600000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
        RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
        RECT 0.74700000 0.18900000 0.79200000 0.20700000 ;
        RECT 1.07100000 0.18900000 1.11600000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.53100000 0.06300000 0.65700000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.14400000 ;
      RECT 0.85500000 0.06300000 0.98100000 0.08100000 ;
      RECT 0.93600000 0.08100000 0.95400000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.85500000 0.18900000 0.98100000 0.20700000 ;
  END

END CKINVDCx8_ASAP7_75t_L
MACRO DFFHQNx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFHQNX1_ASAP7_75T_L 0 0 ;
 SIZE  1.0800000000000007 BY 0.2700000000000002 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.08000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.08000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.01700000 0.06300000 1.06200000 0.08100000 ;
        RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
        RECT 1.01700000 0.18900000 1.06200000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.08300000 ;
      RECT 0.66600000 0.10500000 0.68400000 0.14400000 ;
      RECT 0.93400000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.16400000 ;
      RECT 0.77400000 0.12600000 0.79200000 0.16400000 ;
      RECT 0.01800000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
      RECT 0.55800000 0.06300000 0.60300000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.20900000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.39600000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.39600000 0.20700000 0.41400000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.41400000 0.24300000 ;
      RECT 0.50400000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.50400000 0.22500000 0.54600000 0.24300000 ;
      RECT 0.58900000 0.22500000 0.65700000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.06300000 ;
      RECT 0.80100000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
      RECT 0.85500000 0.02700000 0.90000000 0.04500000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.45000000 0.06300000 0.59600000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.82800000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.77400000 0.14400000 0.90000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.58800000 0.20700000 ;
      RECT 0.51600000 0.22500000 0.61700000 0.24300000 ;
     LAYER V1 ;
      RECT 0.45000000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.57800000 0.06300000 0.59600000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.82800000 0.10700000 0.84600000 0.12500000 ;
      RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.36000000 0.16200000 ;
      RECT 0.45000000 0.14400000 0.46800000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.77400000 0.14400000 0.79200000 0.16200000 ;
      RECT 0.88200000 0.14400000 0.90000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.46600000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.52300000 0.22500000 0.54100000 0.24300000 ;
      RECT 0.59200000 0.22500000 0.61000000 0.24300000 ;
  END

END DFFHQNx1_ASAP7_75t_L
MACRO OA211x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA211X2_ASAP7_75T_L 0 0 ;
 SIZE  0.4320000000000001 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.22500000 ;
        RECT 0.31500000 0.22500000 0.36000000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.17100000 0.04500000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.30600000 0.20700000 ;
      RECT 0.23400000 0.20700000 0.25200000 0.22500000 ;
      RECT 0.18800000 0.22500000 0.25200000 0.24300000 ;
  END

END OA211x2_ASAP7_75t_L
MACRO DFFHQx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFHQX4_ASAP7_75T_L 0 0 ;
 SIZE  1.3500000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.35000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.35000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.12500000 0.06300000 1.25100000 0.08100000 ;
        RECT 1.15200000 0.08100000 1.17000000 0.18900000 ;
        RECT 1.12500000 0.18900000 1.25100000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.63900000 0.02700000 0.71100000 0.04500000 ;
      RECT 0.69300000 0.04500000 0.71100000 0.06300000 ;
      RECT 0.69300000 0.06300000 0.73800000 0.08100000 ;
      RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.08300000 ;
      RECT 0.66600000 0.10500000 0.68400000 0.14400000 ;
      RECT 0.93400000 0.06300000 0.98100000 0.08100000 ;
      RECT 0.96300000 0.08100000 0.98100000 0.10700000 ;
      RECT 0.96300000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.16400000 ;
      RECT 0.09900000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.09900000 0.04500000 0.11700000 0.06300000 ;
      RECT 0.26100000 0.04500000 0.27900000 0.06300000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.26100000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.54800000 0.06300000 0.58600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.55000000 0.18900000 0.58700000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
      RECT 1.01700000 0.06300000 1.06200000 0.08100000 ;
      RECT 1.04400000 0.08100000 1.06200000 0.14500000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.14500000 ;
      RECT 1.04400000 0.14500000 1.11600000 0.16300000 ;
      RECT 1.04400000 0.16300000 1.06200000 0.18900000 ;
      RECT 1.01700000 0.18900000 1.06200000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.39600000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.39600000 0.20700000 0.41400000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.41400000 0.24300000 ;
      RECT 0.50400000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.50400000 0.22500000 0.54100000 0.24300000 ;
      RECT 0.58000000 0.22500000 0.62900000 0.24300000 ;
      RECT 0.81800000 0.06300000 0.85500000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.90000000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.45000000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.71800000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.58500000 0.20700000 ;
      RECT 0.51200000 0.22500000 0.62900000 0.24300000 ;
     LAYER V1 ;
      RECT 0.45000000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.55800000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.71800000 0.06300000 0.73600000 0.08100000 ;
      RECT 0.82800000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.93600000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.36000000 0.16200000 ;
      RECT 0.45000000 0.14400000 0.46800000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.46600000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.51800000 0.22500000 0.53600000 0.24300000 ;
      RECT 0.59600000 0.22500000 0.61400000 0.24300000 ;
  END

END DFFHQx4_ASAP7_75t_L
MACRO OAI333xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI333XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN C3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END C3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.06300000 0.57600000 0.08100000 ;
        RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.57600000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.14400000 ;
    END
  END B3

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
  END

END OAI333xp33_ASAP7_75t_L
MACRO NAND2x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND2X2_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.15300000 0.08100000 0.17100000 0.10700000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.17100000 0.12500000 ;
        RECT 0.28800000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.42300000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.49500000 0.04500000 ;
  END

END NAND2x2_ASAP7_75t_L
MACRO NOR2x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR2X1_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
        RECT 0.18000000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END NOR2x1_ASAP7_75t_L
MACRO AOI31xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI31XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.22500000 0.22500000 0.24300000 ;
  END

END AOI31xp33_ASAP7_75t_L
MACRO NAND2x1p5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND2X1P5_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.12600000 0.11700000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.38700000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
  END

END NAND2x1p5_ASAP7_75t_L
MACRO AOI211x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI211X1_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.12600000 0.11700000 0.16300000 ;
    END
  END A2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
        RECT 0.50400000 0.18900000 0.54900000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.10700000 0.57600000 0.14400000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.36900000 0.22500000 0.60300000 0.24300000 ;
  END

END AOI211x1_ASAP7_75t_L
MACRO NAND2xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND2XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.216 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.21600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.21600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.22500000 ;
        RECT 0.09900000 0.22500000 0.19800000 0.24300000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B

  OBS

  END

END NAND2xp33_ASAP7_75t_L
MACRO OA331x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA331X1_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
        RECT 0.01800000 0.22500000 0.06300000 0.24300000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END B3

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.31500000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.15300000 0.06300000 0.38700000 0.08100000 ;
      RECT 0.47700000 0.06300000 0.52200000 0.08100000 ;
      RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
      RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
      RECT 0.07200000 0.18900000 0.52200000 0.20700000 ;
  END

END OA331x1_ASAP7_75t_L
MACRO ICGx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX2_ASAP7_75T_L 0 0 ;
 SIZE  1.0260000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.02600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.02600000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END SE

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
        RECT 0.61200000 0.10500000 0.63000000 0.18900000 ;
        RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
        RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
       LAYER M2 ;
        RECT 0.34200000 0.10700000 0.63000000 0.12500000 ;
       LAYER V1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
        RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
    END
  END CLK

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.90900000 0.06300000 0.95400000 0.08100000 ;
        RECT 0.93600000 0.08100000 0.95400000 0.22500000 ;
        RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
    END
  END GCLK

  OBS
     LAYER M1 ;
      RECT 0.55600000 0.02700000 0.84600000 0.04500000 ;
      RECT 0.66600000 0.04500000 0.68400000 0.14400000 ;
      RECT 0.82800000 0.04500000 0.84600000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.16500000 ;
      RECT 0.09900000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.28800000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.31500000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.38600000 0.04500000 0.40400000 0.06300000 ;
      RECT 0.38600000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.26100000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.47700000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.47700000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.55800000 0.06300000 0.60300000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.22500000 ;
      RECT 0.55800000 0.22500000 0.60300000 0.24300000 ;
      RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.90000000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
     LAYER M2 ;
      RECT 0.42100000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.35900000 0.18900000 0.57600000 0.20700000 ;
     LAYER V1 ;
      RECT 0.42100000 0.02700000 0.43900000 0.04500000 ;
      RECT 0.55800000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.50400000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.36500000 0.18900000 0.38300000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
  END

END ICGx2_ASAP7_75t_L
MACRO SDFHx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFHX1_ASAP7_75T_L 0 0 ;
 SIZE  1.3500000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.35000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.35000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END D

  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END SI

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.84600000 0.06300000 0.98100000 0.08100000 ;
        RECT 0.28800000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
       LAYER M2 ;
        RECT 0.31300000 0.06300000 0.86600000 0.08100000 ;
       LAYER V1 ;
        RECT 0.31300000 0.06300000 0.33100000 0.08100000 ;
        RECT 0.84800000 0.06300000 0.86600000 0.08100000 ;
    END
  END SE

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.28700000 0.06300000 1.33200000 0.08100000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.22500000 ;
        RECT 1.28700000 0.22500000 1.33200000 0.24300000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.49500000 0.08100000 ;
      RECT 0.82800000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.55800000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.10700000 ;
      RECT 0.50200000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 1.19700000 0.06300000 1.23400000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.14500000 ;
      RECT 0.33200000 0.14500000 0.36900000 0.16300000 ;
      RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.10700000 ;
      RECT 0.18000000 0.10700000 0.25200000 0.12500000 ;
      RECT 0.18000000 0.12500000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.26100000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.82800000 0.14500000 0.89600000 0.16300000 ;
      RECT 0.82800000 0.16300000 0.84600000 0.18900000 ;
      RECT 0.81800000 0.18900000 0.85500000 0.20700000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.18900000 ;
      RECT 1.20400000 0.18900000 1.27800000 0.20700000 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.27900000 0.24300000 ;
      RECT 0.31500000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.68400000 0.20700000 ;
      RECT 0.53100000 0.20700000 0.54900000 0.22500000 ;
      RECT 0.47500000 0.22500000 0.54900000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.73800000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.22500000 ;
      RECT 0.77400000 0.22500000 0.85100000 0.24300000 ;
      RECT 0.85500000 0.02700000 1.03500000 0.04500000 ;
      RECT 1.01700000 0.04500000 1.03500000 0.14500000 ;
      RECT 1.01700000 0.14500000 1.06200000 0.16300000 ;
      RECT 1.01700000 0.16300000 1.03500000 0.18900000 ;
      RECT 0.93600000 0.18900000 1.07200000 0.20700000 ;
      RECT 0.93600000 0.20700000 0.95400000 0.22500000 ;
      RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
      RECT 1.07100000 0.02700000 1.11600000 0.04500000 ;
      RECT 1.09800000 0.04500000 1.11600000 0.22500000 ;
      RECT 1.05000000 0.22500000 1.11600000 0.24300000 ;
      RECT 1.15200000 0.02700000 1.22700000 0.04500000 ;
      RECT 1.15200000 0.04500000 1.17000000 0.22500000 ;
      RECT 1.15200000 0.22500000 1.23100000 0.24300000 ;
     LAYER M2 ;
      RECT 0.96100000 0.06300000 1.22400000 0.08100000 ;
      RECT 0.23200000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 1.17000000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.84600000 0.20700000 ;
      RECT 1.04200000 0.18900000 1.22400000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.49500000 0.24300000 ;
     LAYER V1 ;
      RECT 0.96100000 0.06300000 0.97900000 0.08100000 ;
      RECT 1.20600000 0.06300000 1.22400000 0.08100000 ;
      RECT 0.23200000 0.10700000 0.25000000 0.12500000 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.84800000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 0.36000000 0.16300000 ;
      RECT 1.15200000 0.14500000 1.17000000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.68200000 0.20700000 ;
      RECT 0.82800000 0.18900000 0.84600000 0.20700000 ;
      RECT 1.04200000 0.18900000 1.06000000 0.20700000 ;
      RECT 1.20600000 0.18900000 1.22400000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.27700000 0.24300000 ;
      RECT 0.47700000 0.22500000 0.49500000 0.24300000 ;
  END

END SDFHx1_ASAP7_75t_L
MACRO AOI21xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI21XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.25200000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.25200000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.18900000 0.17100000 0.20700000 ;
  END

END AOI21xp5_ASAP7_75t_L
MACRO AOI22xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI22XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END AOI22xp33_ASAP7_75t_L
MACRO HB4xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HB4XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.31500000 0.18900000 0.36000000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.09000000 0.04500000 ;
      RECT 0.07200000 0.04500000 0.09000000 0.06300000 ;
      RECT 0.07200000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.10700000 ;
      RECT 0.18000000 0.10700000 0.30600000 0.12500000 ;
      RECT 0.28800000 0.12500000 0.30600000 0.14400000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
      RECT 0.04500000 0.22500000 0.09000000 0.24300000 ;
  END

END HB4xp67_ASAP7_75t_L
MACRO AO33x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO33X2_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.22500000 ;
        RECT 0.07200000 0.22500000 0.11700000 0.24300000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B3

  OBS
     LAYER M1 ;
      RECT 0.12600000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.20700000 0.22500000 0.44100000 0.24300000 ;
  END

END AO33x2_ASAP7_75t_L
MACRO ICGx6p67DC_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX6P67DC_ASAP7_75T_L 0 0 ;
 SIZE  2.5920000000000005 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 2.59200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 2.59200000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.09800000 0.12600000 1.11600000 0.16300000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.15200000 0.12600000 1.17000000 0.16300000 ;
    END
  END SE

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.61200000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.22500000 ;
        RECT 0.07200000 0.22500000 1.25100000 0.24300000 ;
        RECT 1.93500000 0.06300000 1.98000000 0.08100000 ;
        RECT 2.47500000 0.06300000 2.52000000 0.08100000 ;
        RECT 1.96200000 0.08100000 1.98000000 0.22500000 ;
        RECT 2.50200000 0.08100000 2.52000000 0.22500000 ;
        RECT 1.55500000 0.22500000 2.52000000 0.24300000 ;
       LAYER M2 ;
        RECT 1.23100000 0.22500000 1.57500000 0.24300000 ;
       LAYER V1 ;
        RECT 1.23100000 0.22500000 1.24900000 0.24300000 ;
        RECT 1.55700000 0.22500000 1.57500000 0.24300000 ;
    END
  END GCLK

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10500000 0.30600000 0.14400000 ;
        RECT 0.82800000 0.10500000 0.84600000 0.14400000 ;
        RECT 0.93600000 0.10500000 0.95400000 0.14400000 ;
        RECT 1.26000000 0.06300000 1.38600000 0.08100000 ;
        RECT 1.26000000 0.08100000 1.27800000 0.14400000 ;
        RECT 1.36800000 0.08100000 1.38600000 0.16400000 ;
       LAYER M2 ;
        RECT 0.28800000 0.10700000 1.27800000 0.12500000 ;
       LAYER V1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.82800000 0.10700000 0.84600000 0.12500000 ;
        RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
        RECT 1.26000000 0.10700000 1.27800000 0.12500000 ;
    END
  END CLK

  OBS
     LAYER M1 ;
      RECT 1.52000000 0.06300000 1.55700000 0.08100000 ;
      RECT 1.53000000 0.08100000 1.54800000 0.12500000 ;
      RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 2.04300000 0.06300000 2.16900000 0.08100000 ;
      RECT 2.12400000 0.08100000 2.14200000 0.14400000 ;
      RECT 1.69200000 0.02700000 2.41200000 0.04500000 ;
      RECT 1.69200000 0.04500000 1.71000000 0.06300000 ;
      RECT 1.63800000 0.06300000 1.71000000 0.08100000 ;
      RECT 1.69200000 0.08100000 1.71000000 0.14400000 ;
      RECT 1.85400000 0.04500000 1.87200000 0.14400000 ;
      RECT 2.23200000 0.04500000 2.25000000 0.14400000 ;
      RECT 2.39400000 0.04500000 2.41200000 0.14400000 ;
      RECT 1.63800000 0.12600000 1.65600000 0.16400000 ;
      RECT 1.80000000 0.12600000 1.81800000 0.16400000 ;
      RECT 2.28600000 0.12600000 2.30400000 0.16400000 ;
      RECT 0.23400000 0.06300000 0.27900000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.54900000 0.20700000 ;
      RECT 0.77400000 0.06300000 0.81900000 0.08100000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.18900000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.66600000 0.18900000 0.87300000 0.20700000 ;
      RECT 0.96300000 0.06300000 1.00800000 0.08100000 ;
      RECT 0.99000000 0.08100000 1.00800000 0.18900000 ;
      RECT 0.95600000 0.18900000 1.00800000 0.20700000 ;
      RECT 1.04400000 0.06300000 1.22400000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
      RECT 1.04400000 0.18900000 1.08900000 0.20700000 ;
      RECT 1.31400000 0.12600000 1.33200000 0.18900000 ;
      RECT 1.12300000 0.18900000 1.38600000 0.20700000 ;
      RECT 1.58400000 0.02700000 1.62900000 0.04500000 ;
      RECT 1.58400000 0.04500000 1.60200000 0.18900000 ;
      RECT 1.55500000 0.18900000 1.62900000 0.20700000 ;
      RECT 1.74600000 0.06300000 1.79100000 0.08100000 ;
      RECT 1.74600000 0.08100000 1.76400000 0.18900000 ;
      RECT 1.90800000 0.12600000 1.92600000 0.18900000 ;
      RECT 1.71900000 0.18900000 1.92600000 0.20700000 ;
      RECT 2.07000000 0.12600000 2.08800000 0.18900000 ;
      RECT 2.04300000 0.18900000 2.16900000 0.20700000 ;
      RECT 2.31300000 0.06300000 2.35800000 0.08100000 ;
      RECT 2.34000000 0.08100000 2.35800000 0.18900000 ;
      RECT 2.44800000 0.12600000 2.46600000 0.18900000 ;
      RECT 2.25900000 0.18900000 2.46600000 0.20700000 ;
      RECT 0.18000000 0.02700000 1.44000000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.14400000 ;
      RECT 0.34200000 0.04500000 0.36000000 0.14400000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.14400000 ;
      RECT 1.42200000 0.04500000 1.44000000 0.22500000 ;
      RECT 1.28700000 0.22500000 1.44000000 0.24300000 ;
      RECT 1.47600000 0.02700000 1.53900000 0.04500000 ;
      RECT 1.47600000 0.04500000 1.49400000 0.22500000 ;
      RECT 1.47600000 0.22500000 1.52100000 0.24300000 ;
     LAYER M2 ;
      RECT 1.53000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14400000 2.30400000 0.16200000 ;
      RECT 0.96300000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.57500000 0.20700000 ;
     LAYER V1 ;
      RECT 1.53000000 0.06300000 1.54800000 0.08100000 ;
      RECT 1.64000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14400000 1.38600000 0.16200000 ;
      RECT 1.63800000 0.14400000 1.65600000 0.16200000 ;
      RECT 1.80000000 0.14400000 1.81800000 0.16200000 ;
      RECT 2.28600000 0.14400000 2.30400000 0.16200000 ;
      RECT 0.96300000 0.18900000 0.98100000 0.20700000 ;
      RECT 1.12500000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.38400000 0.20700000 ;
      RECT 1.55700000 0.18900000 1.57500000 0.20700000 ;
  END

END ICGx6p67DC_ASAP7_75t_L
MACRO AO22x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO22X1_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.06300000 0.30600000 0.08100000 ;
      RECT 0.28800000 0.08100000 0.30600000 0.10700000 ;
      RECT 0.28800000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
      RECT 0.28800000 0.12500000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.30600000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END AO22x1_ASAP7_75t_L
MACRO ICGx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX3_ASAP7_75T_L 0 0 ;
 SIZE  1.0800000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.08000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.08000000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END SE

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
        RECT 0.61200000 0.10500000 0.63000000 0.18900000 ;
        RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
        RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
       LAYER M2 ;
        RECT 0.34200000 0.10700000 0.63000000 0.12500000 ;
       LAYER V1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
        RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
    END
  END CLK

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.90900000 0.06300000 0.95400000 0.08100000 ;
        RECT 0.93600000 0.08100000 0.95400000 0.10700000 ;
        RECT 1.01700000 0.06300000 1.03500000 0.10700000 ;
        RECT 0.93600000 0.10700000 1.03500000 0.12500000 ;
        RECT 1.01700000 0.12500000 1.03500000 0.20700000 ;
        RECT 0.93600000 0.12500000 0.95400000 0.22500000 ;
        RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
    END
  END GCLK

  OBS
     LAYER M1 ;
      RECT 0.55600000 0.02700000 0.84600000 0.04500000 ;
      RECT 0.66600000 0.04500000 0.68400000 0.14400000 ;
      RECT 0.82800000 0.04500000 0.84600000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.16500000 ;
      RECT 0.09900000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.28800000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.31500000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.38600000 0.04500000 0.40400000 0.06300000 ;
      RECT 0.38600000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.26100000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.47700000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.47700000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.55800000 0.06300000 0.60300000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.22500000 ;
      RECT 0.55800000 0.22500000 0.60300000 0.24300000 ;
      RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.90000000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
     LAYER M2 ;
      RECT 0.42100000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.36100000 0.18900000 0.57600000 0.20700000 ;
     LAYER V1 ;
      RECT 0.42100000 0.02700000 0.43900000 0.04500000 ;
      RECT 0.55800000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.50400000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.36600000 0.18900000 0.38400000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
  END

END ICGx3_ASAP7_75t_L
MACRO SDFHx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFHX4_ASAP7_75T_L 0 0 ;
 SIZE  1.6740000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.67400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.67400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END CLK

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.28800000 0.12500000 0.30600000 0.14400000 ;
        RECT 0.54900000 0.10700000 0.58600000 0.12500000 ;
        RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
       LAYER M2 ;
        RECT 0.39400000 0.10700000 0.57600000 0.12500000 ;
       LAYER V1 ;
        RECT 0.39400000 0.10700000 0.41200000 0.12500000 ;
        RECT 0.55800000 0.10700000 0.57600000 0.12500000 ;
    END
  END SE

  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.10700000 0.63000000 0.14400000 ;
    END
  END SI

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.44900000 0.06300000 1.57500000 0.08100000 ;
        RECT 1.47600000 0.08100000 1.49400000 0.18900000 ;
        RECT 1.44900000 0.18900000 1.57500000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.65700000 0.04500000 ;
      RECT 0.69300000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.12700000 ;
      RECT 0.77400000 0.02700000 0.84600000 0.04500000 ;
      RECT 0.82800000 0.04500000 0.84600000 0.08300000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 1.04200000 0.06300000 1.11600000 0.08100000 ;
      RECT 1.09800000 0.08100000 1.11600000 0.14400000 ;
      RECT 0.34000000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.14500000 ;
      RECT 0.65600000 0.14500000 0.69300000 0.16300000 ;
      RECT 0.82800000 0.12600000 0.84600000 0.14500000 ;
      RECT 0.81900000 0.14500000 0.85600000 0.16300000 ;
      RECT 0.04500000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.23400000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.23400000 0.18900000 0.52200000 0.20700000 ;
      RECT 0.58500000 0.18900000 0.76500000 0.20700000 ;
      RECT 0.92700000 0.10700000 0.96400000 0.12500000 ;
      RECT 0.93600000 0.12500000 0.95400000 0.18900000 ;
      RECT 0.80100000 0.18900000 0.95400000 0.20700000 ;
      RECT 1.04400000 0.12600000 1.06200000 0.18900000 ;
      RECT 1.15200000 0.12600000 1.17000000 0.18900000 ;
      RECT 1.04400000 0.18900000 1.17000000 0.20700000 ;
      RECT 1.20600000 0.06300000 1.30500000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.18900000 ;
      RECT 1.20600000 0.18900000 1.30500000 0.20700000 ;
      RECT 0.15300000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.42300000 0.22500000 0.65700000 0.24300000 ;
      RECT 0.99000000 0.02700000 1.08900000 0.04500000 ;
      RECT 0.99000000 0.04500000 1.00800000 0.06300000 ;
      RECT 0.88200000 0.06300000 1.00800000 0.08100000 ;
      RECT 0.88200000 0.08100000 0.90000000 0.14400000 ;
      RECT 0.99000000 0.08100000 1.00800000 0.22500000 ;
      RECT 0.96300000 0.22500000 1.00800000 0.24300000 ;
      RECT 1.12500000 0.02700000 1.35900000 0.04500000 ;
      RECT 1.34100000 0.04500000 1.35900000 0.10700000 ;
      RECT 1.34100000 0.10700000 1.44000000 0.12500000 ;
      RECT 1.42200000 0.12500000 1.44000000 0.14400000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.14500000 ;
      RECT 1.34100000 0.12500000 1.35900000 0.14500000 ;
      RECT 1.26000000 0.14500000 1.35900000 0.16300000 ;
      RECT 1.34100000 0.16300000 1.35900000 0.22500000 ;
      RECT 1.07100000 0.22500000 1.35900000 0.24300000 ;
     LAYER M2 ;
      RECT 0.66400000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.82800000 0.06300000 1.06200000 0.08100000 ;
      RECT 0.72000000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.12600000 0.14500000 0.36000000 0.16300000 ;
      RECT 0.39400000 0.14500000 1.06200000 0.16300000 ;
     LAYER V1 ;
      RECT 0.66400000 0.06300000 0.68200000 0.08100000 ;
      RECT 0.77400000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.82800000 0.06300000 0.84600000 0.08100000 ;
      RECT 1.04400000 0.06300000 1.06200000 0.08100000 ;
      RECT 0.72000000 0.10700000 0.73800000 0.12500000 ;
      RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.12600000 0.14500000 0.14400000 0.16300000 ;
      RECT 0.34200000 0.14500000 0.36000000 0.16300000 ;
      RECT 0.39400000 0.14500000 0.41200000 0.16300000 ;
      RECT 0.66600000 0.14500000 0.68400000 0.16300000 ;
      RECT 0.82800000 0.14500000 0.84600000 0.16300000 ;
      RECT 1.04400000 0.14500000 1.06200000 0.16300000 ;
  END

END SDFHx4_ASAP7_75t_L
MACRO AOI21xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI21XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.25200000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.25200000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.18900000 0.17100000 0.20700000 ;
  END

END AOI21xp33_ASAP7_75t_L
MACRO ICGx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX1_ASAP7_75T_L 0 0 ;
 SIZE  0.9720000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.97200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.97200000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END SE

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
        RECT 0.61200000 0.10500000 0.63000000 0.18900000 ;
        RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
        RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
       LAYER M2 ;
        RECT 0.34200000 0.10700000 0.63000000 0.12500000 ;
       LAYER V1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
        RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
    END
  END CLK

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.90900000 0.06300000 0.95400000 0.08100000 ;
        RECT 0.93600000 0.08100000 0.95400000 0.22500000 ;
        RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
    END
  END GCLK

  OBS
     LAYER M1 ;
      RECT 0.55600000 0.02700000 0.84600000 0.04500000 ;
      RECT 0.66600000 0.04500000 0.68400000 0.14400000 ;
      RECT 0.82800000 0.04500000 0.84600000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.16500000 ;
      RECT 0.09900000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.28800000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.31500000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.38600000 0.04500000 0.40400000 0.06300000 ;
      RECT 0.38600000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.26100000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.47700000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.47700000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.55800000 0.06300000 0.60300000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.22500000 ;
      RECT 0.55800000 0.22500000 0.60300000 0.24300000 ;
      RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.90000000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
     LAYER M2 ;
      RECT 0.42100000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.36100000 0.18900000 0.57600000 0.20700000 ;
     LAYER V1 ;
      RECT 0.42100000 0.02700000 0.43900000 0.04500000 ;
      RECT 0.55800000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.50400000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.36600000 0.18900000 0.38400000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
  END

END ICGx1_ASAP7_75t_L
MACRO INVx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX4_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx4_ASAP7_75t_L
MACRO CKINVDCx5p33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX5P33_ASAP7_75T_L 0 0 ;
 SIZE  1.188 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.18800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.18800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.14500000 ;
        RECT 0.39600000 0.12600000 0.41400000 0.14500000 ;
        RECT 0.72000000 0.12600000 0.73800000 0.14500000 ;
        RECT 1.04400000 0.12600000 1.06200000 0.14500000 ;
        RECT 0.12600000 0.14500000 0.17100000 0.16300000 ;
        RECT 0.36900000 0.14500000 0.41400000 0.16300000 ;
        RECT 0.69300000 0.14500000 0.73800000 0.16300000 ;
        RECT 1.01700000 0.14500000 1.06200000 0.16300000 ;
        RECT 0.15300000 0.16300000 0.17100000 0.22500000 ;
        RECT 0.36900000 0.16300000 0.38700000 0.22500000 ;
        RECT 0.69300000 0.16300000 0.71100000 0.22500000 ;
        RECT 1.01700000 0.16300000 1.03500000 0.22500000 ;
        RECT 0.15300000 0.22500000 1.03500000 0.24300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.02700000 1.03500000 0.04500000 ;
        RECT 0.12600000 0.04500000 0.14400000 0.06300000 ;
        RECT 1.01700000 0.04500000 1.03500000 0.06300000 ;
        RECT 0.07200000 0.06300000 0.14400000 0.08100000 ;
        RECT 1.01700000 0.06300000 1.11600000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.45000000 0.04500000 0.46800000 0.18900000 ;
        RECT 0.77400000 0.04500000 0.79200000 0.18900000 ;
        RECT 1.09800000 0.08100000 1.11600000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
        RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
        RECT 0.74700000 0.18900000 0.79200000 0.20700000 ;
        RECT 1.07100000 0.18900000 1.11600000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.53100000 0.06300000 0.65700000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.14400000 ;
      RECT 0.85500000 0.06300000 0.98100000 0.08100000 ;
      RECT 0.93600000 0.08100000 0.95400000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.85500000 0.18900000 0.98100000 0.20700000 ;
  END

END CKINVDCx5p33_ASAP7_75t_L
MACRO AO31x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO31X2_ASAP7_75T_L 0 0 ;
 SIZE  0.864 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.86400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.86400000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.12600000 0.11700000 0.16300000 ;
    END
  END A3

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
        RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
        RECT 0.74700000 0.18900000 0.79200000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.36900000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
      RECT 0.31500000 0.04500000 0.33300000 0.06300000 ;
      RECT 0.31500000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.20700000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.53100000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.14500000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.14500000 ;
      RECT 0.55800000 0.14500000 0.73800000 0.16300000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.55800000 0.16300000 0.57600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.54900000 0.24300000 ;
  END

END AO31x2_ASAP7_75t_L
MACRO OA33x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA33X2_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.22500000 ;
        RECT 0.07200000 0.22500000 0.11700000 0.24300000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A3

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B1

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.12600000 0.06300000 0.49500000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.33300000 0.20700000 ;
  END

END OA33x2_ASAP7_75t_L
MACRO NOR4xp75_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR4XP75_ASAP7_75T_L 0 0 ;
 SIZE  0.756 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.75600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.75600000 0.27900000 ;
    END
  END VDD

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END D

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
        RECT 0.58500000 0.18900000 0.71100000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.66600000 0.12600000 0.68400000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.09900000 0.22500000 0.33300000 0.24300000 ;
      RECT 0.42300000 0.22500000 0.65700000 0.24300000 ;
  END

END NOR4xp75_ASAP7_75t_L
MACRO DECAPx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DECAPX2_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  OBS
     LAYER M1 ;
      RECT 0.12600000 0.06300000 0.27900000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.18000000 0.12600000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
  END

END DECAPx2_ASAP7_75t_L
MACRO OA31x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA31X2_ASAP7_75T_L 0 0 ;
 SIZE  0.81 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.81000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.81000000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.12600000 0.22500000 0.16300000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.12600000 0.44100000 0.16300000 ;
    END
  END A3

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END B1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.69300000 0.06300000 0.73800000 0.08100000 ;
        RECT 0.72000000 0.08100000 0.73800000 0.18900000 ;
        RECT 0.69300000 0.18900000 0.73800000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.04500000 0.18900000 0.27900000 0.20700000 ;
      RECT 0.04500000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.14500000 ;
      RECT 0.61200000 0.14500000 0.68400000 0.16300000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
      RECT 0.61200000 0.16300000 0.63000000 0.18900000 ;
      RECT 0.34200000 0.18900000 0.63000000 0.20700000 ;
      RECT 0.20700000 0.22500000 0.44100000 0.24300000 ;
  END

END OA31x2_ASAP7_75t_L
MACRO NOR3x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR3X2_ASAP7_75T_L 0 0 ;
 SIZE  1.08 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.08000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.08000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.02700000 0.95400000 0.04500000 ;
        RECT 0.18000000 0.04500000 0.19800000 0.06300000 ;
        RECT 0.12600000 0.06300000 0.19800000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.93600000 0.04500000 0.95400000 0.18900000 ;
        RECT 0.04500000 0.18900000 0.17100000 0.20700000 ;
        RECT 0.90900000 0.18900000 1.03500000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.06300000 0.90000000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.10700000 ;
        RECT 0.18000000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.18000000 0.12500000 0.19800000 0.14400000 ;
        RECT 0.88200000 0.08100000 0.90000000 0.14400000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.14500000 ;
        RECT 0.72000000 0.12600000 0.73800000 0.14500000 ;
        RECT 0.34200000 0.14500000 0.49500000 0.16300000 ;
        RECT 0.58500000 0.14500000 0.73800000 0.16300000 ;
        RECT 0.47700000 0.16300000 0.49500000 0.18900000 ;
        RECT 0.58500000 0.16300000 0.60300000 0.18900000 ;
        RECT 0.47700000 0.18900000 0.60300000 0.20700000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.53100000 0.12600000 0.54900000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.22500000 0.33300000 0.24300000 ;
      RECT 0.26100000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.66600000 0.18900000 0.81900000 0.20700000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.66600000 0.20700000 0.68400000 0.22500000 ;
      RECT 0.42300000 0.22500000 0.68400000 0.24300000 ;
      RECT 0.74700000 0.22500000 0.98100000 0.24300000 ;
  END

END NOR3x2_ASAP7_75t_L
MACRO XNOR2x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XNOR2X1_ASAP7_75T_L 0 0 ;
 SIZE  0.6480000000000001 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
        RECT 0.44800000 0.10700000 0.52200000 0.12500000 ;
        RECT 0.50400000 0.12500000 0.52200000 0.14400000 ;
       LAYER M2 ;
        RECT 0.34200000 0.10700000 0.46800000 0.12500000 ;
       LAYER V1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
        RECT 0.45000000 0.10700000 0.46800000 0.12500000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.28800000 0.12500000 0.30600000 0.18900000 ;
        RECT 0.55800000 0.12600000 0.57600000 0.18900000 ;
        RECT 0.28800000 0.18900000 0.57600000 0.20700000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.06300000 0.63000000 0.08100000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.63000000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.16400000 ;
      RECT 0.01800000 0.02700000 0.17100000 0.04500000 ;
      RECT 0.20700000 0.14400000 0.25200000 0.16200000 ;
      RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
      RECT 0.20700000 0.16200000 0.22500000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.22500000 0.20700000 ;
     LAYER M2 ;
      RECT 0.23200000 0.14400000 0.41400000 0.16200000 ;
     LAYER V1 ;
      RECT 0.23200000 0.14400000 0.25000000 0.16200000 ;
      RECT 0.39600000 0.14400000 0.41400000 0.16200000 ;
  END

END XNOR2x1_ASAP7_75t_L
MACRO OAI22x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI22X1_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.22500000 ;
        RECT 0.04500000 0.22500000 0.52200000 0.24300000 ;
    END
  END Y

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.14500000 ;
        RECT 0.07200000 0.14500000 0.11700000 0.16300000 ;
        RECT 0.09900000 0.16300000 0.11700000 0.18900000 ;
        RECT 0.23400000 0.12600000 0.25200000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.25200000 0.20700000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.14500000 ;
        RECT 0.42300000 0.14500000 0.46800000 0.16300000 ;
        RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
        RECT 0.42300000 0.16300000 0.44100000 0.18900000 ;
        RECT 0.28800000 0.18900000 0.44100000 0.20700000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.36900000 0.12600000 0.38700000 0.16300000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.49500000 0.04500000 ;
  END

END OAI22x1_ASAP7_75t_L
MACRO DFFHQNx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFHQNX2_ASAP7_75T_L 0 0 ;
 SIZE  1.0260000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.02600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.02600000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.85500000 0.06300000 0.90000000 0.08100000 ;
        RECT 0.88200000 0.08100000 0.90000000 0.22500000 ;
        RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.61200000 0.06300000 0.66200000 0.08100000 ;
      RECT 0.64400000 0.08100000 0.66200000 0.10700000 ;
      RECT 0.60600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.23400000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.61000000 0.14700000 0.68400000 0.16500000 ;
      RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.18000000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.45000000 0.14500000 0.46800000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.42300000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.55800000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.55800000 0.04500000 0.57600000 0.22500000 ;
      RECT 0.55800000 0.22500000 0.60300000 0.24300000 ;
      RECT 0.69300000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.18900000 ;
      RECT 0.82800000 0.12600000 0.84600000 0.18900000 ;
      RECT 0.66600000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.66600000 0.20700000 0.68400000 0.22500000 ;
      RECT 0.63900000 0.22500000 0.68400000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.98100000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 0.93600000 0.04500000 0.95400000 0.22500000 ;
      RECT 0.93600000 0.22500000 0.98100000 0.24300000 ;
     LAYER M2 ;
      RECT 0.44800000 0.06300000 0.63200000 0.08100000 ;
      RECT 0.12600000 0.10700000 0.25200000 0.12500000 ;
      RECT 0.45000000 0.14700000 0.63000000 0.16500000 ;
     LAYER V1 ;
      RECT 0.44800000 0.06300000 0.46600000 0.08100000 ;
      RECT 0.61400000 0.06300000 0.63200000 0.08100000 ;
      RECT 0.12600000 0.10700000 0.14400000 0.12500000 ;
      RECT 0.23400000 0.10700000 0.25200000 0.12500000 ;
      RECT 0.45000000 0.14700000 0.46800000 0.16500000 ;
      RECT 0.61200000 0.14700000 0.63000000 0.16500000 ;
  END

END DFFHQNx2_ASAP7_75t_L
MACRO O2A1O1Ixp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN O2A1O1IXP5_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.25200000 0.08100000 ;
        RECT 0.09900000 0.08100000 0.11700000 0.10700000 ;
        RECT 0.07200000 0.10700000 0.11700000 0.12500000 ;
        RECT 0.07200000 0.12500000 0.09000000 0.14400000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.36900000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.15300000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.09900000 0.22500000 0.22500000 0.24300000 ;
  END

END O2A1O1Ixp5_ASAP7_75t_L
MACRO OR3x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR3X1_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.30600000 0.04500000 ;
        RECT 0.28800000 0.04500000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
  END

END OR3x1_ASAP7_75t_L
MACRO CKINVDCx11_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX11_ASAP7_75T_L 0 0 ;
 SIZE  1.4040000000000001 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.40400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.40400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.38700000 0.04500000 ;
        RECT 0.15300000 0.04500000 0.17100000 0.10700000 ;
        RECT 0.36900000 0.04500000 0.38700000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.17100000 0.12500000 ;
        RECT 0.36900000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
        RECT 0.85500000 0.06300000 0.98100000 0.08100000 ;
        RECT 1.28700000 0.06300000 1.33200000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.22500000 ;
        RECT 0.88200000 0.08100000 0.90000000 0.22500000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.22500000 ;
        RECT 0.07200000 0.22500000 1.33200000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.63900000 0.06300000 0.76500000 0.08100000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 0.58500000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.58500000 0.04500000 0.60300000 0.10700000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.10700000 ;
      RECT 0.55800000 0.10700000 0.60300000 0.12500000 ;
      RECT 0.80100000 0.10700000 0.84600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.82800000 0.12500000 0.84600000 0.14400000 ;
      RECT 1.07100000 0.06300000 1.19700000 0.08100000 ;
      RECT 1.15200000 0.08100000 1.17000000 0.14400000 ;
      RECT 1.01700000 0.02700000 1.25100000 0.04500000 ;
      RECT 1.01700000 0.04500000 1.03500000 0.10700000 ;
      RECT 1.23300000 0.04500000 1.25100000 0.10700000 ;
      RECT 0.99000000 0.10700000 1.03500000 0.12500000 ;
      RECT 1.23300000 0.10700000 1.27800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 1.26000000 0.12500000 1.27800000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.63900000 0.18900000 0.76500000 0.20700000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.18900000 ;
      RECT 1.07100000 0.18900000 1.19700000 0.20700000 ;
  END

END CKINVDCx11_ASAP7_75t_L
MACRO AND5x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND5X1_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END D

  PIN E
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END E

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.36900000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.22500000 ;
        RECT 0.36900000 0.22500000 0.41400000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.36000000 0.20700000 ;
  END

END AND5x1_ASAP7_75t_L
MACRO AOI332xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI332XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
        RECT 0.42300000 0.18900000 0.52200000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.26100000 0.22500000 0.49500000 0.24300000 ;
  END

END AOI332xp33_ASAP7_75t_L
MACRO A2O1A1O1Ixp25_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN A2O1A1O1IXP25_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.38700000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.34200000 0.18900000 0.44100000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END D

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.04500000 0.22500000 0.17100000 0.24300000 ;
      RECT 0.20700000 0.22500000 0.38700000 0.24300000 ;
  END

END A2O1A1O1Ixp25_ASAP7_75t_L
MACRO HB3xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HB3XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.09000000 0.04500000 ;
      RECT 0.07200000 0.04500000 0.09000000 0.06300000 ;
      RECT 0.07200000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.10700000 ;
      RECT 0.18000000 0.10700000 0.25200000 0.12500000 ;
      RECT 0.23400000 0.12500000 0.25200000 0.14400000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
      RECT 0.04500000 0.22500000 0.09000000 0.24300000 ;
  END

END HB3xp67_ASAP7_75t_L
MACRO ICGx2p67DC_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX2P67DC_ASAP7_75T_L 0 0 ;
 SIZE  2.5920000000000005 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 2.59200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 2.59200000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.09800000 0.12600000 1.11600000 0.16300000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.15200000 0.12600000 1.17000000 0.16300000 ;
    END
  END SE

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.61200000 0.02700000 0.65700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.22500000 ;
        RECT 0.61200000 0.04500000 0.63000000 0.22500000 ;
        RECT 0.07200000 0.22500000 1.25100000 0.24300000 ;
        RECT 1.93500000 0.02700000 1.98000000 0.04500000 ;
        RECT 2.47500000 0.02700000 2.52000000 0.04500000 ;
        RECT 1.96200000 0.04500000 1.98000000 0.22500000 ;
        RECT 2.50200000 0.04500000 2.52000000 0.22500000 ;
        RECT 1.55500000 0.22500000 2.52000000 0.24300000 ;
       LAYER M2 ;
        RECT 1.23100000 0.22500000 1.57500000 0.24300000 ;
       LAYER V1 ;
        RECT 1.23100000 0.22500000 1.24900000 0.24300000 ;
        RECT 1.55700000 0.22500000 1.57500000 0.24300000 ;
    END
  END GCLK

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10500000 0.30600000 0.14400000 ;
        RECT 0.82800000 0.10500000 0.84600000 0.14400000 ;
        RECT 0.93600000 0.10500000 0.95400000 0.14400000 ;
        RECT 1.26000000 0.06300000 1.38600000 0.08100000 ;
        RECT 1.26000000 0.08100000 1.27800000 0.14400000 ;
        RECT 1.36800000 0.08100000 1.38600000 0.14500000 ;
        RECT 1.35900000 0.14500000 1.39500000 0.16300000 ;
       LAYER M2 ;
        RECT 0.28800000 0.10700000 1.27800000 0.12500000 ;
       LAYER V1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.82800000 0.10700000 0.84600000 0.12500000 ;
        RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
        RECT 1.26000000 0.10700000 1.27800000 0.12500000 ;
    END
  END CLK

  OBS
     LAYER M1 ;
      RECT 1.52000000 0.06300000 1.55700000 0.08100000 ;
      RECT 1.53000000 0.08100000 1.54800000 0.12500000 ;
      RECT 0.18000000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.14400000 ;
      RECT 0.34200000 0.04500000 0.36000000 0.14400000 ;
      RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 1.71900000 0.02700000 1.89900000 0.04500000 ;
      RECT 1.71900000 0.04500000 1.73700000 0.06300000 ;
      RECT 1.63800000 0.06300000 1.73700000 0.08100000 ;
      RECT 1.69200000 0.08100000 1.71000000 0.14400000 ;
      RECT 1.85400000 0.04500000 1.87200000 0.14400000 ;
      RECT 2.04300000 0.06300000 2.19600000 0.08100000 ;
      RECT 2.17800000 0.08100000 2.19600000 0.14400000 ;
      RECT 2.01400000 0.02700000 2.41200000 0.04500000 ;
      RECT 2.23200000 0.04500000 2.25000000 0.14400000 ;
      RECT 2.39400000 0.04500000 2.41200000 0.14400000 ;
      RECT 1.74600000 0.12600000 1.76400000 0.14500000 ;
      RECT 1.74000000 0.14500000 1.77000000 0.16300000 ;
      RECT 2.06800000 0.14500000 2.14200000 0.16300000 ;
      RECT 2.28600000 0.12600000 2.30400000 0.14500000 ;
      RECT 2.28000000 0.14500000 2.31000000 0.16300000 ;
      RECT 1.63800000 0.12600000 1.65600000 0.16500000 ;
      RECT 0.23400000 0.06300000 0.27900000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.54900000 0.20700000 ;
      RECT 0.77400000 0.06300000 0.81900000 0.08100000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.18900000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.66600000 0.18900000 0.87300000 0.20700000 ;
      RECT 0.96300000 0.06300000 1.00800000 0.08100000 ;
      RECT 0.99000000 0.08100000 1.00800000 0.18900000 ;
      RECT 0.95800000 0.18900000 1.00800000 0.20700000 ;
      RECT 1.04400000 0.06300000 1.22400000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
      RECT 1.04400000 0.18900000 1.08900000 0.20700000 ;
      RECT 1.31400000 0.12600000 1.33200000 0.18900000 ;
      RECT 1.12300000 0.18900000 1.38800000 0.20700000 ;
      RECT 1.58400000 0.02700000 1.62900000 0.04500000 ;
      RECT 1.58400000 0.04500000 1.60200000 0.18900000 ;
      RECT 1.53000000 0.18900000 1.62900000 0.20700000 ;
      RECT 1.77300000 0.06300000 1.81800000 0.08100000 ;
      RECT 1.80000000 0.08100000 1.81800000 0.18900000 ;
      RECT 1.90800000 0.12600000 1.92600000 0.18900000 ;
      RECT 1.71900000 0.18900000 1.92600000 0.20700000 ;
      RECT 2.01600000 0.12600000 2.03400000 0.18900000 ;
      RECT 2.01600000 0.18900000 2.16900000 0.20700000 ;
      RECT 2.31300000 0.06300000 2.35800000 0.08100000 ;
      RECT 2.34000000 0.08100000 2.35800000 0.18900000 ;
      RECT 2.44800000 0.12700000 2.46600000 0.18900000 ;
      RECT 2.25900000 0.18900000 2.46600000 0.20700000 ;
      RECT 0.69100000 0.02700000 1.44000000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.14400000 ;
      RECT 1.42200000 0.04500000 1.44000000 0.22500000 ;
      RECT 1.28700000 0.22500000 1.44000000 0.24300000 ;
      RECT 1.47600000 0.02700000 1.54100000 0.04500000 ;
      RECT 1.47600000 0.04500000 1.49400000 0.22500000 ;
      RECT 1.47600000 0.22500000 1.52100000 0.24300000 ;
     LAYER M2 ;
      RECT 0.55600000 0.02700000 0.71100000 0.04500000 ;
      RECT 1.87900000 0.02700000 2.03400000 0.04500000 ;
      RECT 1.53000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14500000 2.08800000 0.16300000 ;
      RECT 2.12200000 0.14500000 2.30400000 0.16300000 ;
      RECT 0.96300000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36800000 0.18900000 1.55200000 0.20700000 ;
     LAYER V1 ;
      RECT 0.55600000 0.02700000 0.57400000 0.04500000 ;
      RECT 0.69300000 0.02700000 0.71100000 0.04500000 ;
      RECT 1.87900000 0.02700000 1.89700000 0.04500000 ;
      RECT 2.01600000 0.02700000 2.03400000 0.04500000 ;
      RECT 1.53000000 0.06300000 1.54800000 0.08100000 ;
      RECT 1.64000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14500000 1.38600000 0.16300000 ;
      RECT 1.63800000 0.14500000 1.65600000 0.16300000 ;
      RECT 1.74600000 0.14500000 1.76400000 0.16300000 ;
      RECT 2.07000000 0.14500000 2.08800000 0.16300000 ;
      RECT 2.12200000 0.14500000 2.14000000 0.16300000 ;
      RECT 2.28600000 0.14500000 2.30400000 0.16300000 ;
      RECT 0.96300000 0.18900000 0.98100000 0.20700000 ;
      RECT 1.12500000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36800000 0.18900000 1.38600000 0.20700000 ;
      RECT 1.53400000 0.18900000 1.55200000 0.20700000 ;
  END

END ICGx2p67DC_ASAP7_75t_L
MACRO AOI321xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI321XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.31500000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.22500000 0.22500000 0.24300000 ;
      RECT 0.26100000 0.22500000 0.38700000 0.24300000 ;
  END

END AOI321xp33_ASAP7_75t_L
MACRO INVx5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX5_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx5_ASAP7_75t_L
MACRO AOI221x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI221X1_ASAP7_75T_L 0 0 ;
 SIZE  0.756 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.75600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.75600000 0.27900000 ;
    END
  END VDD

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.63000000 0.08100000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
        RECT 0.61200000 0.18900000 0.65700000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B2

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.66600000 0.12600000 0.68400000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.31500000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.04500000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.31500000 0.22500000 0.71100000 0.24300000 ;
  END

END AOI221x1_ASAP7_75t_L
MACRO NOR2x1p5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR2X1P5_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.38700000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.22500000 0.33300000 0.24300000 ;
  END

END NOR2x1p5_ASAP7_75t_L
MACRO OAI22xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI22XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.17100000 0.20700000 ;
    END
  END Y

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END B1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
  END

END OAI22xp33_ASAP7_75t_L
MACRO AND4x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND4X1_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END D

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.22500000 ;
        RECT 0.31500000 0.22500000 0.36000000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.30600000 0.20700000 ;
  END

END AND4x1_ASAP7_75t_L
MACRO OAI22xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI22XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.17100000 0.20700000 ;
    END
  END Y

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END B1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
  END

END OAI22xp5_ASAP7_75t_L
MACRO INVxp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVXP67_ASAP7_75T_L 0 0 ;
 SIZE  0.162 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.16200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.16200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  OBS

  END

END INVxp67_ASAP7_75t_L
MACRO SDFLx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFLX2_ASAP7_75T_L 0 0 ;
 SIZE  1.4040000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.40400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.40400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END D

  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END SI

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16500000 ;
        RECT 1.20600000 0.12600000 1.22400000 0.16500000 ;
       LAYER M2 ;
        RECT 0.28800000 0.14500000 1.22400000 0.16300000 ;
       LAYER V1 ;
        RECT 0.28800000 0.14500000 0.30600000 0.16300000 ;
        RECT 1.20600000 0.14500000 1.22400000 0.16300000 ;
    END
  END SE

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.28700000 0.06300000 1.33200000 0.08100000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.18900000 ;
        RECT 1.28700000 0.18900000 1.33200000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.42300000 0.06300000 0.60300000 0.08100000 ;
      RECT 0.85300000 0.10700000 0.90000000 0.12500000 ;
      RECT 0.34200000 0.06100000 0.36000000 0.14400000 ;
      RECT 0.61200000 0.10500000 0.63000000 0.14400000 ;
      RECT 1.26000000 0.10500000 1.27800000 0.14400000 ;
      RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.31500000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.55800000 0.12600000 0.57600000 0.18900000 ;
      RECT 0.66600000 0.14500000 0.68400000 0.18900000 ;
      RECT 0.52900000 0.18900000 0.68400000 0.20700000 ;
      RECT 1.09600000 0.06300000 1.19700000 0.08100000 ;
      RECT 1.15200000 0.08100000 1.17000000 0.18900000 ;
      RECT 1.15200000 0.18900000 1.19700000 0.20700000 ;
      RECT 0.82800000 0.14500000 0.84600000 0.20900000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.26100000 0.22500000 0.49500000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.73800000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.22500000 ;
      RECT 0.77400000 0.22500000 0.81900000 0.24300000 ;
      RECT 0.85500000 0.02700000 0.92700000 0.04500000 ;
      RECT 0.90900000 0.04500000 0.92700000 0.06300000 ;
      RECT 0.90900000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.93600000 0.08100000 0.95400000 0.10700000 ;
      RECT 0.93600000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.93600000 0.12500000 0.95400000 0.22500000 ;
      RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
      RECT 1.04400000 0.02700000 1.08900000 0.04500000 ;
      RECT 1.04400000 0.04500000 1.06200000 0.22500000 ;
      RECT 1.04400000 0.22500000 1.08900000 0.24300000 ;
     LAYER M2 ;
      RECT 0.34200000 0.06300000 1.11600000 0.08100000 ;
      RECT 0.18000000 0.10700000 0.87300000 0.12500000 ;
      RECT 0.98800000 0.10700000 1.27800000 0.12500000 ;
      RECT 0.09900000 0.18900000 0.54900000 0.20700000 ;
      RECT 0.63900000 0.18900000 0.84600000 0.20700000 ;
     LAYER V1 ;
      RECT 0.34200000 0.06300000 0.36000000 0.08100000 ;
      RECT 1.09800000 0.06300000 1.11600000 0.08100000 ;
      RECT 0.18000000 0.10700000 0.19800000 0.12500000 ;
      RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
      RECT 0.85500000 0.10700000 0.87300000 0.12500000 ;
      RECT 0.98800000 0.10700000 1.00600000 0.12500000 ;
      RECT 1.26000000 0.10700000 1.27800000 0.12500000 ;
      RECT 0.09900000 0.18900000 0.11700000 0.20700000 ;
      RECT 0.53100000 0.18900000 0.54900000 0.20700000 ;
      RECT 0.63900000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.82800000 0.18900000 0.84600000 0.20700000 ;
  END

END SDFLx2_ASAP7_75t_L
MACRO DFFASRHQNx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFASRHQNX1_ASAP7_75T_L 0 0 ;
 SIZE  1.4040000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.40400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.40400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN RESETN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.10500000 0.63000000 0.14400000 ;
        RECT 1.04400000 0.10500000 1.06200000 0.14400000 ;
       LAYER M2 ;
        RECT 0.61200000 0.10700000 1.06200000 0.12500000 ;
       LAYER V1 ;
        RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
        RECT 1.04400000 0.10700000 1.06200000 0.12500000 ;
    END
  END RESETN

  PIN SETN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.66600000 0.12600000 0.68400000 0.16400000 ;
        RECT 0.77400000 0.12600000 0.79200000 0.16400000 ;
        RECT 0.99000000 0.12600000 1.00800000 0.16400000 ;
       LAYER M2 ;
        RECT 0.66600000 0.14400000 1.00800000 0.16200000 ;
       LAYER V1 ;
        RECT 0.66600000 0.14400000 0.68400000 0.16200000 ;
        RECT 0.77400000 0.14400000 0.79200000 0.16200000 ;
        RECT 0.99000000 0.14400000 1.00800000 0.16200000 ;
    END
  END SETN

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.34100000 0.06300000 1.38600000 0.08100000 ;
        RECT 1.36800000 0.08100000 1.38600000 0.18900000 ;
        RECT 1.34100000 0.18900000 1.38600000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.39600000 0.06300000 0.43400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.45000000 0.10500000 0.46800000 0.14400000 ;
      RECT 0.69100000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.06300000 ;
      RECT 0.80100000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.14400000 ;
      RECT 0.87200000 0.06300000 0.91000000 0.08100000 ;
      RECT 0.88200000 0.08100000 0.90000000 0.14400000 ;
      RECT 0.93600000 0.06300000 1.03500000 0.08100000 ;
      RECT 0.93600000 0.08100000 0.95400000 0.14400000 ;
      RECT 0.85500000 0.02700000 1.27800000 0.04500000 ;
      RECT 1.26000000 0.04500000 1.27800000 0.10700000 ;
      RECT 1.26000000 0.10700000 1.33200000 0.12500000 ;
      RECT 1.31400000 0.12500000 1.33200000 0.14400000 ;
      RECT 1.26000000 0.12500000 1.27800000 0.16400000 ;
      RECT 0.15300000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.34200000 0.04500000 0.36000000 0.14400000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.42300000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.18900000 ;
      RECT 0.36900000 0.18900000 0.52200000 0.20700000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.69100000 0.18900000 0.73800000 0.20700000 ;
      RECT 0.77400000 0.18900000 0.81900000 0.20700000 ;
      RECT 0.23400000 0.06300000 0.30600000 0.08100000 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.25200000 0.24300000 ;
      RECT 0.42300000 0.22500000 0.60300000 0.24300000 ;
      RECT 0.58500000 0.02700000 0.65700000 0.04500000 ;
      RECT 0.58500000 0.04500000 0.60300000 0.06300000 ;
      RECT 0.63900000 0.04500000 0.65700000 0.06300000 ;
      RECT 0.55800000 0.06300000 0.60300000 0.08100000 ;
      RECT 0.63900000 0.06300000 0.76500000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.55800000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.63900000 0.20700000 0.65700000 0.22500000 ;
      RECT 0.63900000 0.22500000 0.81900000 0.24300000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.18900000 ;
      RECT 0.88200000 0.18900000 1.11600000 0.20700000 ;
      RECT 0.88200000 0.20700000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
      RECT 0.93400000 0.22500000 0.98100000 0.24300000 ;
      RECT 1.07100000 0.22500000 1.11600000 0.24300000 ;
      RECT 1.15200000 0.18700000 1.17000000 0.22500000 ;
      RECT 1.15200000 0.22500000 1.19700000 0.24300000 ;
      RECT 1.06900000 0.06300000 1.17000000 0.08100000 ;
      RECT 1.15200000 0.08100000 1.17000000 0.10700000 ;
      RECT 1.15200000 0.10700000 1.22400000 0.12500000 ;
      RECT 1.15200000 0.12500000 1.17000000 0.14400000 ;
      RECT 1.20600000 0.12500000 1.22400000 0.18900000 ;
      RECT 1.20600000 0.18900000 1.28700000 0.20700000 ;
      RECT 1.26900000 0.20700000 1.28700000 0.22500000 ;
      RECT 1.23100000 0.22500000 1.28700000 0.24300000 ;
     LAYER M2 ;
      RECT 0.36700000 0.02700000 0.71100000 0.04500000 ;
      RECT 0.28600000 0.06300000 0.90000000 0.08100000 ;
      RECT 1.01500000 0.06300000 1.08900000 0.08100000 ;
      RECT 0.34200000 0.10700000 0.46800000 0.12500000 ;
      RECT 1.09800000 0.14400000 1.27800000 0.16200000 ;
      RECT 0.47700000 0.18900000 0.71100000 0.20700000 ;
      RECT 0.79900000 0.18900000 1.17000000 0.20700000 ;
      RECT 0.79900000 0.22500000 0.95400000 0.24300000 ;
      RECT 1.09600000 0.22500000 1.25100000 0.24300000 ;
     LAYER V1 ;
      RECT 0.36700000 0.02700000 0.38500000 0.04500000 ;
      RECT 0.69300000 0.02700000 0.71100000 0.04500000 ;
      RECT 0.28600000 0.06300000 0.30400000 0.08100000 ;
      RECT 0.41100000 0.06300000 0.42900000 0.08100000 ;
      RECT 0.88200000 0.06300000 0.90000000 0.08100000 ;
      RECT 1.01500000 0.06300000 1.03300000 0.08100000 ;
      RECT 1.07100000 0.06300000 1.08900000 0.08100000 ;
      RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
      RECT 0.45000000 0.10700000 0.46800000 0.12500000 ;
      RECT 1.09800000 0.14400000 1.11600000 0.16200000 ;
      RECT 1.26000000 0.14400000 1.27800000 0.16200000 ;
      RECT 0.47700000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.69300000 0.18900000 0.71100000 0.20700000 ;
      RECT 0.79900000 0.18900000 0.81700000 0.20700000 ;
      RECT 1.15200000 0.18900000 1.17000000 0.20700000 ;
      RECT 0.79900000 0.22500000 0.81700000 0.24300000 ;
      RECT 0.93600000 0.22500000 0.95400000 0.24300000 ;
      RECT 1.09600000 0.22500000 1.11400000 0.24300000 ;
      RECT 1.23300000 0.22500000 1.25100000 0.24300000 ;
  END

END DFFASRHQNx1_ASAP7_75t_L
MACRO AOI33xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI33XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A3

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.22500000 0.33300000 0.24300000 ;
  END

END AOI33xp33_ASAP7_75t_L
MACRO OR4x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR4X2_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.18900000 ;
        RECT 0.18000000 0.18900000 0.22500000 0.20700000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.06300000 0.27900000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
        RECT 0.28800000 0.18900000 0.33300000 0.20700000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.18000000 0.02700000 0.41400000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.06300000 ;
      RECT 0.12600000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.39600000 0.04500000 0.41400000 0.18900000 ;
      RECT 0.36900000 0.18900000 0.41400000 0.20700000 ;
  END

END OR4x2_ASAP7_75t_L
MACRO OAI331xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI331XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
      RECT 0.26100000 0.06300000 0.38700000 0.08100000 ;
  END

END OAI331xp33_ASAP7_75t_L
MACRO CKINVDCx14_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX14_ASAP7_75T_L 0 0 ;
 SIZE  1.512 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.51200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.51200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.38700000 0.04500000 ;
        RECT 0.15300000 0.04500000 0.17100000 0.10700000 ;
        RECT 0.36900000 0.04500000 0.38700000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.17100000 0.12500000 ;
        RECT 0.36900000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.85500000 0.02700000 1.27800000 0.04500000 ;
        RECT 1.26000000 0.04500000 1.27800000 0.06300000 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
        RECT 1.26000000 0.06300000 1.41300000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.93600000 0.04500000 0.95400000 0.18900000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.14400000 0.20700000 ;
        RECT 0.80100000 0.18900000 0.98100000 0.20700000 ;
        RECT 1.28700000 0.18900000 1.41300000 0.20700000 ;
        RECT 0.12600000 0.20700000 0.14400000 0.22500000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.22500000 ;
        RECT 0.80100000 0.20700000 0.81900000 0.22500000 ;
        RECT 0.12600000 0.22500000 0.81900000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.63900000 0.06300000 0.76500000 0.08100000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 0.58500000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.58500000 0.04500000 0.60300000 0.10700000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.10700000 ;
      RECT 0.55800000 0.10700000 0.60300000 0.12500000 ;
      RECT 0.80100000 0.10700000 0.84600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.82800000 0.12500000 0.84600000 0.14400000 ;
      RECT 1.07100000 0.06300000 1.19700000 0.08100000 ;
      RECT 1.15200000 0.08100000 1.17000000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.63900000 0.18900000 0.76500000 0.20700000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.18900000 ;
      RECT 1.07100000 0.18900000 1.19700000 0.20700000 ;
      RECT 0.99000000 0.12600000 1.00800000 0.14500000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.14500000 ;
      RECT 0.99000000 0.14500000 1.03500000 0.16300000 ;
      RECT 1.23300000 0.14500000 1.27800000 0.16300000 ;
      RECT 1.01700000 0.16300000 1.03500000 0.22500000 ;
      RECT 1.23300000 0.16300000 1.25100000 0.22500000 ;
      RECT 1.01700000 0.22500000 1.25100000 0.24300000 ;
  END

END CKINVDCx14_ASAP7_75t_L
MACRO DHLx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DHLX1_ASAP7_75T_L 0 0 ;
 SIZE  0.8100000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.81000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.81000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
        RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
        RECT 0.74700000 0.18900000 0.79200000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.50400000 0.10500000 0.52200000 0.14400000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.14500000 ;
      RECT 0.66400000 0.14500000 0.73800000 0.16300000 ;
      RECT 0.07200000 0.02700000 0.33300000 0.04500000 ;
      RECT 0.07200000 0.04500000 0.09000000 0.06300000 ;
      RECT 0.31500000 0.04500000 0.33300000 0.06300000 ;
      RECT 0.01800000 0.06300000 0.09000000 0.08100000 ;
      RECT 0.31500000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.41400000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.42300000 0.02700000 0.54900000 0.04500000 ;
      RECT 0.53100000 0.04500000 0.54900000 0.06300000 ;
      RECT 0.53100000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.50400000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.50400000 0.20700000 0.52200000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.58500000 0.02700000 0.63000000 0.04500000 ;
      RECT 0.61200000 0.04500000 0.63000000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.63000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.50400000 0.10700000 0.63000000 0.12500000 ;
      RECT 0.55800000 0.14500000 0.68400000 0.16300000 ;
     LAYER V1 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
      RECT 0.55800000 0.14500000 0.57600000 0.16300000 ;
      RECT 0.66600000 0.14500000 0.68400000 0.16300000 ;
  END

END DHLx1_ASAP7_75t_L
MACRO OA222x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA222X2_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END C1

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.53100000 0.06300000 0.57600000 0.08100000 ;
        RECT 0.55800000 0.08100000 0.57600000 0.22500000 ;
        RECT 0.53100000 0.22500000 0.57600000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.20700000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.52200000 0.20700000 ;
  END

END OA222x2_ASAP7_75t_L
MACRO ICGx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX4_ASAP7_75T_L 0 0 ;
 SIZE  1.1340000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.13400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.13400000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END SE

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
        RECT 0.61200000 0.10500000 0.63000000 0.18900000 ;
        RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
        RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
       LAYER M2 ;
        RECT 0.34200000 0.10700000 0.63000000 0.12500000 ;
       LAYER V1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.12500000 ;
        RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
    END
  END CLK

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.90900000 0.06300000 1.03500000 0.08100000 ;
        RECT 0.93600000 0.08100000 0.95400000 0.18900000 ;
        RECT 0.93600000 0.18900000 1.03500000 0.20700000 ;
        RECT 0.93600000 0.20700000 0.95400000 0.22500000 ;
        RECT 0.90900000 0.22500000 0.95400000 0.24300000 ;
    END
  END GCLK

  OBS
     LAYER M1 ;
      RECT 0.55600000 0.02700000 0.84600000 0.04500000 ;
      RECT 0.66600000 0.04500000 0.68400000 0.14400000 ;
      RECT 0.82800000 0.04500000 0.84600000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.16500000 ;
      RECT 0.09900000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.28800000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.31500000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.38600000 0.04500000 0.40400000 0.06300000 ;
      RECT 0.38600000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.26100000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.47700000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.47700000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.55800000 0.06300000 0.60300000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.22500000 ;
      RECT 0.55800000 0.22500000 0.60300000 0.24300000 ;
      RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.90000000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
     LAYER M2 ;
      RECT 0.42100000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.36100000 0.18900000 0.57600000 0.20700000 ;
     LAYER V1 ;
      RECT 0.42100000 0.02700000 0.43900000 0.04500000 ;
      RECT 0.55800000 0.02700000 0.57600000 0.04500000 ;
      RECT 0.39600000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.50400000 0.14500000 0.52200000 0.16300000 ;
      RECT 0.36600000 0.18900000 0.38400000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
  END

END ICGx4_ASAP7_75t_L
MACRO NOR3x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR3X1_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.42300000 0.18900000 0.54900000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.26100000 0.22500000 0.49500000 0.24300000 ;
  END

END NOR3x1_ASAP7_75t_L
MACRO CKINVDCx16_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX16_ASAP7_75T_L 0 0 ;
 SIZE  1.62 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.62000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.62000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.49500000 0.04500000 ;
        RECT 0.26100000 0.04500000 0.27900000 0.10700000 ;
        RECT 0.47700000 0.04500000 0.49500000 0.10700000 ;
        RECT 0.23400000 0.10700000 0.27900000 0.12500000 ;
        RECT 0.47700000 0.10700000 0.52200000 0.12500000 ;
        RECT 0.23400000 0.12500000 0.25200000 0.14400000 ;
        RECT 0.50400000 0.12500000 0.52200000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.96300000 0.02700000 1.52100000 0.04500000 ;
        RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.53100000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
        RECT 1.04400000 0.04500000 1.06200000 0.18900000 ;
        RECT 1.42200000 0.04500000 1.44000000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.19800000 0.20700000 ;
        RECT 1.04400000 0.18900000 1.08900000 0.20700000 ;
        RECT 1.39500000 0.18900000 1.52100000 0.20700000 ;
        RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
        RECT 0.55800000 0.08100000 0.57600000 0.22500000 ;
        RECT 1.04400000 0.20700000 1.06200000 0.22500000 ;
        RECT 0.18000000 0.22500000 1.06200000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.31500000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.74700000 0.06300000 0.87300000 0.08100000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.14400000 ;
      RECT 0.69300000 0.02700000 0.92700000 0.04500000 ;
      RECT 0.69300000 0.04500000 0.71100000 0.10700000 ;
      RECT 0.90900000 0.04500000 0.92700000 0.10700000 ;
      RECT 0.66600000 0.10700000 0.71100000 0.12500000 ;
      RECT 0.90900000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.66600000 0.12500000 0.68400000 0.14400000 ;
      RECT 0.93600000 0.12500000 0.95400000 0.14400000 ;
      RECT 1.17900000 0.06300000 1.30500000 0.08100000 ;
      RECT 1.26000000 0.08100000 1.27800000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
      RECT 0.31500000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.82800000 0.12600000 0.84600000 0.18900000 ;
      RECT 0.74700000 0.18900000 0.87300000 0.20700000 ;
      RECT 1.20600000 0.12600000 1.22400000 0.18900000 ;
      RECT 1.17900000 0.18900000 1.30500000 0.20700000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.14500000 ;
      RECT 1.36800000 0.12600000 1.38600000 0.14500000 ;
      RECT 1.09800000 0.14500000 1.14300000 0.16300000 ;
      RECT 1.34100000 0.14500000 1.38600000 0.16300000 ;
      RECT 1.12500000 0.16300000 1.14300000 0.22500000 ;
      RECT 1.34100000 0.16300000 1.35900000 0.22500000 ;
      RECT 1.12500000 0.22500000 1.35900000 0.24300000 ;
  END

END CKINVDCx16_ASAP7_75t_L
MACRO OAI332xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI332XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.52200000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.14400000 ;
    END
  END B3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
  END

END OAI332xp33_ASAP7_75t_L
MACRO DFFLQNx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFLQNX2_ASAP7_75T_L 0 0 ;
 SIZE  1.1340000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.13400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.13400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.01700000 0.06300000 1.06200000 0.08100000 ;
        RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
        RECT 1.01700000 0.18900000 1.06200000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.08300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.08300000 ;
      RECT 0.66600000 0.10500000 0.68400000 0.14400000 ;
      RECT 0.93400000 0.06300000 0.98100000 0.08100000 ;
      RECT 0.96300000 0.08100000 0.98100000 0.10700000 ;
      RECT 0.96300000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.16400000 ;
      RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.06300000 ;
      RECT 0.18000000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
      RECT 0.54800000 0.06300000 0.58500000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.20900000 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.28800000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
      RECT 0.28800000 0.20700000 0.30600000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.30600000 0.24300000 ;
      RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.50400000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.50400000 0.22500000 0.54100000 0.24300000 ;
      RECT 0.59000000 0.22500000 0.65700000 0.24300000 ;
      RECT 0.81800000 0.06300000 0.85600000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.90000000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.45000000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.72000000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.58200000 0.20700000 ;
      RECT 0.51400000 0.22500000 0.61900000 0.24300000 ;
     LAYER V1 ;
      RECT 0.45000000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.55800000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.72000000 0.06300000 0.73800000 0.08100000 ;
      RECT 0.82800000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.93600000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.36000000 0.16200000 ;
      RECT 0.45000000 0.14400000 0.46800000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.46600000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.52100000 0.22500000 0.53900000 0.24300000 ;
      RECT 0.59400000 0.22500000 0.61200000 0.24300000 ;
  END

END DFFLQNx2_ASAP7_75t_L
MACRO AND4x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND4X2_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.07200000 0.22500000 0.11700000 0.24300000 ;
    END
  END Y

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.36900000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.41400000 0.20700000 ;
  END

END AND4x2_ASAP7_75t_L
MACRO NAND5xp2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND5XP2_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.27900000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END D

  PIN E
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END E

  OBS

  END

END NAND5xp2_ASAP7_75t_L
MACRO OR2x6_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR2X6_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
        RECT 0.09900000 0.20700000 0.11700000 0.22500000 ;
        RECT 0.23400000 0.12600000 0.25200000 0.22500000 ;
        RECT 0.09900000 0.22500000 0.25200000 0.24300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.02700000 0.36000000 0.04500000 ;
        RECT 0.34200000 0.04500000 0.36000000 0.06300000 ;
        RECT 0.34200000 0.06300000 0.54900000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.31500000 0.18900000 0.54900000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.30600000 0.08100000 ;
      RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
  END

END OR2x6_ASAP7_75t_L
MACRO SDFLx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFLX1_ASAP7_75T_L 0 0 ;
 SIZE  1.3500000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.35000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.35000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END D

  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END SI

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.84600000 0.06300000 0.95400000 0.08100000 ;
        RECT 0.28800000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
       LAYER M2 ;
        RECT 0.31300000 0.06300000 0.86600000 0.08100000 ;
       LAYER V1 ;
        RECT 0.31300000 0.06300000 0.33100000 0.08100000 ;
        RECT 0.84800000 0.06300000 0.86600000 0.08100000 ;
    END
  END SE

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.28700000 0.06300000 1.33200000 0.08100000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.22500000 ;
        RECT 1.28700000 0.22500000 1.33200000 0.24300000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.49500000 0.08100000 ;
      RECT 0.81900000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.55800000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.10700000 ;
      RECT 0.50200000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 1.17700000 0.06300000 1.22400000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.14500000 ;
      RECT 0.33300000 0.14500000 0.37000000 0.16300000 ;
      RECT 0.04500000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.10700000 ;
      RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
      RECT 0.12600000 0.12500000 0.14400000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.26100000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.82800000 0.14500000 0.90200000 0.16300000 ;
      RECT 0.82800000 0.16300000 0.84600000 0.18900000 ;
      RECT 0.81900000 0.18900000 0.85900000 0.20700000 ;
      RECT 1.12500000 0.02700000 1.19700000 0.04500000 ;
      RECT 1.12500000 0.04500000 1.14300000 0.14500000 ;
      RECT 1.09600000 0.14500000 1.17000000 0.16300000 ;
      RECT 1.15200000 0.16300000 1.17000000 0.18900000 ;
      RECT 1.15200000 0.18900000 1.19700000 0.20700000 ;
      RECT 0.15300000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.20700000 0.04500000 0.22500000 0.06300000 ;
      RECT 0.20700000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14500000 ;
      RECT 0.20700000 0.14500000 0.25200000 0.16300000 ;
      RECT 0.20700000 0.16300000 0.22500000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.27900000 0.24300000 ;
      RECT 0.31500000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.68400000 0.20700000 ;
      RECT 0.53100000 0.20700000 0.54900000 0.22500000 ;
      RECT 0.47500000 0.22500000 0.54900000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.73800000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.22500000 ;
      RECT 0.77400000 0.22500000 0.85900000 0.24300000 ;
      RECT 0.85500000 0.02700000 1.00800000 0.04500000 ;
      RECT 0.99000000 0.04500000 1.00800000 0.18900000 ;
      RECT 0.94900000 0.18900000 1.00800000 0.20700000 ;
      RECT 0.94900000 0.20700000 0.96700000 0.22500000 ;
      RECT 0.90900000 0.22500000 1.00800000 0.24300000 ;
      RECT 1.04400000 0.02700000 1.08900000 0.04500000 ;
      RECT 1.04400000 0.04500000 1.06200000 0.22500000 ;
      RECT 1.04400000 0.22500000 1.08900000 0.24300000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.18900000 ;
      RECT 1.23300000 0.18900000 1.27800000 0.20700000 ;
      RECT 1.23300000 0.20700000 1.25100000 0.22500000 ;
      RECT 1.12300000 0.22500000 1.25100000 0.24300000 ;
     LAYER M2 ;
      RECT 0.93400000 0.06300000 1.19700000 0.08100000 ;
      RECT 0.17800000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 1.11600000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.49500000 0.24300000 ;
      RECT 0.98800000 0.22500000 1.14300000 0.24300000 ;
     LAYER V1 ;
      RECT 0.93400000 0.06300000 0.95200000 0.08100000 ;
      RECT 1.17900000 0.06300000 1.19700000 0.08100000 ;
      RECT 0.17800000 0.10700000 0.19600000 0.12500000 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.84800000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 0.36000000 0.16300000 ;
      RECT 1.09800000 0.14500000 1.11600000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.68200000 0.20700000 ;
      RECT 0.82800000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.27700000 0.24300000 ;
      RECT 0.47700000 0.22500000 0.49500000 0.24300000 ;
      RECT 0.98800000 0.22500000 1.00600000 0.24300000 ;
      RECT 1.12500000 0.22500000 1.14300000 0.24300000 ;
  END

END SDFLx1_ASAP7_75t_L
MACRO SDFLx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFLX3_ASAP7_75T_L 0 0 ;
 SIZE  1.4580000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.45800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.45800000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END D

  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END SI

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.84600000 0.06300000 0.98100000 0.08100000 ;
        RECT 0.28800000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
       LAYER M2 ;
        RECT 0.31300000 0.06300000 0.86600000 0.08100000 ;
       LAYER V1 ;
        RECT 0.31300000 0.06300000 0.33100000 0.08100000 ;
        RECT 0.84800000 0.06300000 0.86600000 0.08100000 ;
    END
  END SE

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.28700000 0.06300000 1.41300000 0.08100000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.18900000 ;
        RECT 1.31400000 0.18900000 1.41300000 0.20700000 ;
        RECT 1.31400000 0.20700000 1.33200000 0.22500000 ;
        RECT 1.28700000 0.22500000 1.33200000 0.24300000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.36900000 0.06300000 0.49500000 0.08100000 ;
      RECT 0.82800000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.55800000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.10700000 ;
      RECT 0.50200000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 1.19600000 0.06300000 1.23700000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.14500000 ;
      RECT 0.33300000 0.14500000 0.37000000 0.16300000 ;
      RECT 0.04500000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.10700000 ;
      RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
      RECT 0.12600000 0.12500000 0.14400000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.26100000 0.18900000 0.49500000 0.20700000 ;
      RECT 0.82800000 0.14500000 0.90000000 0.16300000 ;
      RECT 0.82800000 0.16300000 0.84600000 0.18900000 ;
      RECT 0.81800000 0.18900000 0.85800000 0.20700000 ;
      RECT 1.15200000 0.02700000 1.22400000 0.04500000 ;
      RECT 1.15200000 0.04500000 1.17000000 0.18900000 ;
      RECT 1.15200000 0.18900000 1.19700000 0.20700000 ;
      RECT 0.15300000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.20700000 0.04500000 0.22500000 0.06300000 ;
      RECT 0.20700000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14500000 ;
      RECT 0.20700000 0.14500000 0.25200000 0.16300000 ;
      RECT 0.20700000 0.16300000 0.22500000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.27900000 0.24300000 ;
      RECT 0.31500000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.68400000 0.20700000 ;
      RECT 0.53100000 0.20700000 0.54900000 0.22500000 ;
      RECT 0.47500000 0.22500000 0.54900000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.73800000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.22500000 ;
      RECT 0.77400000 0.22500000 0.85600000 0.24300000 ;
      RECT 0.85500000 0.02700000 1.03500000 0.04500000 ;
      RECT 1.01700000 0.04500000 1.03500000 0.10700000 ;
      RECT 0.99000000 0.10700000 1.06200000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.22500000 ;
      RECT 0.90900000 0.22500000 1.03500000 0.24300000 ;
      RECT 1.07100000 0.02700000 1.11600000 0.04500000 ;
      RECT 1.09800000 0.04500000 1.11600000 0.14500000 ;
      RECT 1.04400000 0.14500000 1.11600000 0.16300000 ;
      RECT 1.09800000 0.16300000 1.11600000 0.22500000 ;
      RECT 1.07100000 0.22500000 1.11600000 0.24300000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.18900000 ;
      RECT 1.23300000 0.18900000 1.27800000 0.20700000 ;
      RECT 1.23300000 0.20700000 1.25100000 0.22500000 ;
      RECT 1.15000000 0.22500000 1.25100000 0.24300000 ;
     LAYER M2 ;
      RECT 0.96100000 0.06300000 1.22400000 0.08100000 ;
      RECT 0.17800000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 1.17000000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.49500000 0.24300000 ;
      RECT 1.01500000 0.22500000 1.17000000 0.24300000 ;
     LAYER V1 ;
      RECT 0.96100000 0.06300000 0.97900000 0.08100000 ;
      RECT 1.20600000 0.06300000 1.22400000 0.08100000 ;
      RECT 0.17800000 0.10700000 0.19600000 0.12500000 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.84800000 0.10700000 0.86600000 0.12500000 ;
      RECT 0.34200000 0.14500000 0.36000000 0.16300000 ;
      RECT 1.15200000 0.14500000 1.17000000 0.16300000 ;
      RECT 0.66400000 0.18900000 0.68200000 0.20700000 ;
      RECT 0.82800000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.25900000 0.22500000 0.27700000 0.24300000 ;
      RECT 0.47700000 0.22500000 0.49500000 0.24300000 ;
      RECT 1.01500000 0.22500000 1.03300000 0.24300000 ;
      RECT 1.15200000 0.22500000 1.17000000 0.24300000 ;
  END

END SDFLx3_ASAP7_75t_L
MACRO BUFx12_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX12_ASAP7_75T_L 0 0 ;
 SIZE  0.864 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.86400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.86400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.76500000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.76500000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.10700000 ;
      RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
      RECT 0.18000000 0.12500000 0.19800000 0.14400000 ;
      RECT 0.12600000 0.12500000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx12_ASAP7_75t_L
MACRO NAND2x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND2X1_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
  END

END NAND2x1_ASAP7_75t_L
MACRO AO331x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO331X1_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.02700000 0.06300000 0.04500000 ;
        RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B3

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.31500000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.07200000 0.06300000 0.52200000 0.08100000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
      RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
      RECT 0.47700000 0.18900000 0.52200000 0.20700000 ;
      RECT 0.15300000 0.22500000 0.38700000 0.24300000 ;
  END

END AO331x1_ASAP7_75t_L
MACRO AO32x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO32X2_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  OBS
     LAYER M1 ;
      RECT 0.12600000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
      RECT 0.36900000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.20700000 0.22500000 0.44100000 0.24300000 ;
  END

END AO32x2_ASAP7_75t_L
MACRO AND3x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND3X2_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.30600000 0.24300000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.23400000 0.12600000 0.25200000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.25200000 0.20700000 ;
  END

END AND3x2_ASAP7_75t_L
MACRO AO322x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO322X2_ASAP7_75T_L 0 0 ;
 SIZE  0.81 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.81000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.81000000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C1

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END C2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.63900000 0.06300000 0.76500000 0.08100000 ;
        RECT 0.72000000 0.08100000 0.73800000 0.18900000 ;
        RECT 0.63900000 0.18900000 0.76500000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.04500000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.14500000 ;
      RECT 0.55800000 0.14500000 0.68400000 0.16300000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
      RECT 0.55800000 0.16300000 0.57600000 0.18900000 ;
      RECT 0.39600000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.26100000 0.22500000 0.49500000 0.24300000 ;
  END

END AO322x2_ASAP7_75t_L
MACRO OAI21x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI21X1_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
        RECT 0.36900000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.22500000 ;
        RECT 0.01800000 0.22500000 0.41400000 0.24300000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
        RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.36000000 0.20700000 ;
    END
  END B

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
  END

END OAI21x1_ASAP7_75t_L
MACRO INVx6_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX6_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx6_ASAP7_75t_L
MACRO OA21x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA21X2_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.30600000 0.04500000 ;
        RECT 0.28800000 0.04500000 0.30600000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.30600000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.17100000 0.04500000 ;
      RECT 0.09900000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.25200000 0.20700000 ;
  END

END OA21x2_ASAP7_75t_L
MACRO BUFx8_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX8_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.54900000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.54900000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.10700000 ;
      RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
      RECT 0.18000000 0.12500000 0.19800000 0.14400000 ;
      RECT 0.12600000 0.12500000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx8_ASAP7_75t_L
MACRO SDFHx2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFHX2_ASAP7_75T_L 0 0 ;
 SIZE  1.4040000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.15200000 0.10700000 1.17000000 0.14400000 ;
    END
  END SI

  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.40400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.40400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.17100000 0.20700000 ;
    END
  END QN

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.82800000 0.12600000 0.84600000 0.16300000 ;
    END
  END D

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.09800000 0.10700000 1.11600000 0.14400000 ;
        RECT 1.20600000 0.10700000 1.22400000 0.14500000 ;
        RECT 1.31400000 0.12600000 1.33200000 0.14500000 ;
        RECT 1.20600000 0.14500000 1.33200000 0.16300000 ;
       LAYER M2 ;
        RECT 1.09800000 0.10900000 1.22400000 0.12700000 ;
       LAYER V1 ;
        RECT 1.09800000 0.10900000 1.11600000 0.12700000 ;
        RECT 1.20600000 0.10900000 1.22400000 0.12700000 ;
    END
  END SE

  OBS
     LAYER M1 ;
      RECT 0.90900000 0.06300000 0.98100000 0.08100000 ;
      RECT 1.01500000 0.06300000 1.19700000 0.08100000 ;
      RECT 0.85500000 0.02700000 0.98100000 0.04500000 ;
      RECT 0.85500000 0.04500000 0.87300000 0.08300000 ;
      RECT 0.45000000 0.10600000 0.46800000 0.14400000 ;
      RECT 0.61200000 0.10500000 0.63000000 0.14400000 ;
      RECT 0.77400000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 0.99000000 0.10500000 1.00800000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.14500000 ;
      RECT 0.28600000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.55800000 0.12600000 0.57600000 0.16500000 ;
      RECT 0.93600000 0.12600000 0.95400000 0.16500000 ;
      RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
      RECT 0.36900000 0.06300000 0.52200000 0.08100000 ;
      RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
      RECT 0.36900000 0.18900000 0.52200000 0.20700000 ;
      RECT 0.63700000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.18900000 ;
      RECT 0.63700000 0.18900000 0.68400000 0.20700000 ;
      RECT 0.95500000 0.18900000 0.99200000 0.20700000 ;
      RECT 1.12300000 0.18900000 1.19700000 0.20700000 ;
      RECT 1.07100000 0.18400000 1.08900000 0.23000000 ;
      RECT 0.19400000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.19400000 0.04500000 0.21200000 0.22500000 ;
      RECT 0.19400000 0.22500000 0.27900000 0.24300000 ;
      RECT 0.31500000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.31500000 0.04500000 0.33300000 0.06300000 ;
      RECT 0.26100000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.26100000 0.08100000 0.27900000 0.10700000 ;
      RECT 0.23400000 0.10700000 0.27900000 0.12500000 ;
      RECT 0.23400000 0.12500000 0.25200000 0.18900000 ;
      RECT 0.23400000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.31500000 0.20700000 0.33300000 0.22500000 ;
      RECT 0.31500000 0.22500000 0.54900000 0.24300000 ;
      RECT 0.80100000 0.22500000 0.87300000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 1.04400000 0.12600000 1.06200000 0.15100000 ;
      RECT 1.01700000 0.15100000 1.06200000 0.16900000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.18800000 ;
      RECT 0.88200000 0.12600000 0.90000000 0.18800000 ;
      RECT 0.72000000 0.18800000 0.92700000 0.20600000 ;
      RECT 0.72000000 0.20600000 0.73800000 0.22500000 ;
      RECT 0.90900000 0.20600000 0.92700000 0.22500000 ;
      RECT 1.01700000 0.16900000 1.03500000 0.22500000 ;
      RECT 0.63900000 0.22500000 0.73800000 0.24300000 ;
      RECT 0.90900000 0.22500000 1.03500000 0.24300000 ;
      RECT 1.11200000 0.22500000 1.20200000 0.24300000 ;
      RECT 1.01500000 0.02700000 1.35900000 0.04500000 ;
      RECT 1.34100000 0.04500000 1.35900000 0.06300000 ;
      RECT 1.34100000 0.06300000 1.38600000 0.08100000 ;
      RECT 1.36800000 0.08100000 1.38600000 0.22500000 ;
      RECT 1.28700000 0.22500000 1.38600000 0.24300000 ;
     LAYER M2 ;
      RECT 0.79900000 0.02700000 1.03500000 0.04500000 ;
      RECT 0.64200000 0.06300000 0.87300000 0.08100000 ;
      RECT 0.96100000 0.06300000 1.03500000 0.08100000 ;
      RECT 0.50400000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.19400000 0.10800000 0.46800000 0.12600000 ;
      RECT 0.01800000 0.14500000 0.30600000 0.16300000 ;
      RECT 0.36900000 0.14500000 0.95400000 0.16300000 ;
      RECT 0.63900000 0.18900000 0.98300000 0.20700000 ;
      RECT 1.07100000 0.18900000 1.14300000 0.20700000 ;
      RECT 0.85300000 0.22500000 1.20000000 0.24300000 ;
     LAYER V1 ;
      RECT 0.79900000 0.02700000 0.81700000 0.04500000 ;
      RECT 1.01700000 0.02700000 1.03500000 0.04500000 ;
      RECT 0.64200000 0.06300000 0.66000000 0.08100000 ;
      RECT 0.85500000 0.06300000 0.87300000 0.08100000 ;
      RECT 0.96100000 0.06300000 0.97900000 0.08100000 ;
      RECT 1.01700000 0.06300000 1.03500000 0.08100000 ;
      RECT 0.50400000 0.10700000 0.52200000 0.12500000 ;
      RECT 0.61200000 0.10700000 0.63000000 0.12500000 ;
      RECT 0.99000000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.19400000 0.10800000 0.21200000 0.12600000 ;
      RECT 0.45000000 0.10800000 0.46800000 0.12600000 ;
      RECT 0.01800000 0.14500000 0.03600000 0.16300000 ;
      RECT 0.28800000 0.14500000 0.30600000 0.16300000 ;
      RECT 0.36900000 0.14500000 0.38700000 0.16300000 ;
      RECT 0.55800000 0.14500000 0.57600000 0.16300000 ;
      RECT 0.93600000 0.14500000 0.95400000 0.16300000 ;
      RECT 0.63900000 0.18900000 0.65700000 0.20700000 ;
      RECT 0.96500000 0.18900000 0.98300000 0.20700000 ;
      RECT 1.07100000 0.18900000 1.08900000 0.20700000 ;
      RECT 1.12500000 0.18900000 1.14300000 0.20700000 ;
      RECT 0.85300000 0.22500000 0.87100000 0.24300000 ;
      RECT 1.18200000 0.22500000 1.20000000 0.24300000 ;
  END

END SDFHx2_ASAP7_75t_L
MACRO BUFx12f_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX12F_ASAP7_75T_L 0 0 ;
 SIZE  0.972 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.97200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.97200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.12600000 0.17100000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.87300000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.31500000 0.18900000 0.87300000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14500000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.14500000 ;
      RECT 0.23400000 0.14500000 0.30600000 0.16300000 ;
      RECT 0.23400000 0.16300000 0.25200000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.25200000 0.20700000 ;
  END

END BUFx12f_ASAP7_75t_L
MACRO NAND4xp25_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND4XP25_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.04500000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END A

  OBS

  END

END NAND4xp25_ASAP7_75t_L
MACRO BUFx4f_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX4F_ASAP7_75T_L 0 0 ;
 SIZE  0.4320000000000001 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.10700000 ;
      RECT 0.12600000 0.10700000 0.19800000 0.12500000 ;
      RECT 0.18000000 0.12500000 0.19800000 0.14400000 ;
      RECT 0.12600000 0.12500000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx4f_ASAP7_75t_L
MACRO BUFx24_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX24_ASAP7_75T_L 0 0 ;
 SIZE  1.62 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.62000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.62000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 1.52100000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.31500000 0.18900000 1.52100000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
      RECT 0.15300000 0.08100000 0.17100000 0.14500000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.14500000 ;
      RECT 0.15300000 0.14500000 0.30600000 0.16300000 ;
      RECT 0.15300000 0.16300000 0.17100000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.17100000 0.20700000 ;
      RECT 0.20700000 0.16300000 0.22500000 0.20700000 ;
  END

END BUFx24_ASAP7_75t_L
MACRO SDFLx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN SDFLX4_ASAP7_75T_L 0 0 ;
 SIZE  1.6740000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.67400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.67400000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END CLK

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.28800000 0.12500000 0.30600000 0.14400000 ;
        RECT 0.54800000 0.10700000 0.58500000 0.12500000 ;
        RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
       LAYER M2 ;
        RECT 0.39400000 0.10700000 0.57600000 0.12500000 ;
       LAYER V1 ;
        RECT 0.39400000 0.10700000 0.41200000 0.12500000 ;
        RECT 0.55800000 0.10700000 0.57600000 0.12500000 ;
    END
  END SE

  PIN SI
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.12600000 0.63000000 0.16300000 ;
    END
  END SI

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.44900000 0.06300000 1.57500000 0.08100000 ;
        RECT 1.47600000 0.08100000 1.49400000 0.18900000 ;
        RECT 1.44900000 0.18900000 1.57500000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.65700000 0.04500000 ;
      RECT 0.69300000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.12700000 ;
      RECT 0.77400000 0.02700000 0.84600000 0.04500000 ;
      RECT 0.82800000 0.04500000 0.84600000 0.08300000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 1.04200000 0.06300000 1.11600000 0.08100000 ;
      RECT 1.09800000 0.08100000 1.11600000 0.14400000 ;
      RECT 0.34000000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.14500000 ;
      RECT 0.65600000 0.14500000 0.69300000 0.16300000 ;
      RECT 0.82800000 0.12600000 0.84600000 0.14500000 ;
      RECT 0.81800000 0.14500000 0.85500000 0.16300000 ;
      RECT 0.09900000 0.02700000 0.38700000 0.04500000 ;
      RECT 0.09900000 0.04500000 0.11700000 0.06300000 ;
      RECT 0.36900000 0.04500000 0.38700000 0.06300000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.36900000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.23400000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.23400000 0.18900000 0.52200000 0.20700000 ;
      RECT 0.58500000 0.18900000 0.76500000 0.20700000 ;
      RECT 0.92700000 0.10700000 0.96400000 0.12500000 ;
      RECT 0.93600000 0.12500000 0.95400000 0.18900000 ;
      RECT 0.80100000 0.18900000 0.95400000 0.20700000 ;
      RECT 1.04400000 0.12600000 1.06200000 0.18900000 ;
      RECT 1.15200000 0.12600000 1.17000000 0.18900000 ;
      RECT 1.04400000 0.18900000 1.17000000 0.20700000 ;
      RECT 1.20600000 0.06300000 1.30500000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.18900000 ;
      RECT 1.20600000 0.18900000 1.30500000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.42300000 0.22500000 0.65700000 0.24300000 ;
      RECT 0.99000000 0.02700000 1.08900000 0.04500000 ;
      RECT 0.99000000 0.04500000 1.00800000 0.06300000 ;
      RECT 0.88200000 0.06300000 1.00800000 0.08100000 ;
      RECT 0.88200000 0.08100000 0.90000000 0.14400000 ;
      RECT 0.99000000 0.08100000 1.00800000 0.22500000 ;
      RECT 0.96300000 0.22500000 1.00800000 0.24300000 ;
      RECT 1.12500000 0.02700000 1.35900000 0.04500000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.14500000 ;
      RECT 1.34100000 0.04500000 1.35900000 0.14500000 ;
      RECT 1.42200000 0.12600000 1.44000000 0.14500000 ;
      RECT 1.26000000 0.14500000 1.44000000 0.16300000 ;
      RECT 1.34100000 0.16300000 1.35900000 0.22500000 ;
      RECT 1.07100000 0.22500000 1.35900000 0.24300000 ;
     LAYER M2 ;
      RECT 0.66400000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.82800000 0.06300000 1.06200000 0.08100000 ;
      RECT 0.72000000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.18000000 0.14500000 0.36000000 0.16300000 ;
      RECT 0.39400000 0.14500000 1.06200000 0.16300000 ;
     LAYER V1 ;
      RECT 0.66400000 0.06300000 0.68200000 0.08100000 ;
      RECT 0.77400000 0.06300000 0.79200000 0.08100000 ;
      RECT 0.82800000 0.06300000 0.84600000 0.08100000 ;
      RECT 1.04400000 0.06300000 1.06200000 0.08100000 ;
      RECT 0.72000000 0.10700000 0.73800000 0.12500000 ;
      RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.18000000 0.14500000 0.19800000 0.16300000 ;
      RECT 0.34200000 0.14500000 0.36000000 0.16300000 ;
      RECT 0.39400000 0.14500000 0.41200000 0.16300000 ;
      RECT 0.66600000 0.14500000 0.68400000 0.16300000 ;
      RECT 0.82800000 0.14500000 0.84600000 0.16300000 ;
      RECT 1.04400000 0.14500000 1.06200000 0.16300000 ;
  END

END SDFLx4_ASAP7_75t_L
MACRO INVx11_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX11_ASAP7_75T_L 0 0 ;
 SIZE  0.7020000000000001 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.70200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.70200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.31500000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.65700000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx11_ASAP7_75t_L
MACRO OAI211xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI211XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.17100000 0.04500000 ;
  END

END OAI211xp5_ASAP7_75t_L
MACRO OR3x4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR3X4_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
        RECT 0.28800000 0.04500000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.38700000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
  END

END OR3x4_ASAP7_75t_L
MACRO HAxp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HAXP5_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
        RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.36000000 0.20700000 ;
    END
  END A

  PIN CON
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
        RECT 0.01800000 0.22500000 0.11700000 0.24300000 ;
    END
  END CON

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.14500000 ;
        RECT 0.28800000 0.12600000 0.30600000 0.14500000 ;
        RECT 0.12600000 0.14500000 0.30600000 0.16300000 ;
    END
  END B

  PIN SN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
        RECT 0.45000000 0.04500000 0.46800000 0.18900000 ;
        RECT 0.39600000 0.18900000 0.46800000 0.20700000 ;
        RECT 0.39600000 0.20700000 0.41400000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.41400000 0.24300000 ;
    END
  END SN

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
  END

END HAxp5_ASAP7_75t_L
MACRO NAND2xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND2XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.32400000000000007 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.06300000 0.22500000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.14500000 ;
        RECT 0.15300000 0.14500000 0.19800000 0.16300000 ;
        RECT 0.15300000 0.16300000 0.17100000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.12600000 0.11700000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
  END

END NAND2xp67_ASAP7_75t_L
MACRO AO21x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO21X1_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.30600000 0.04500000 ;
        RECT 0.28800000 0.04500000 0.30600000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.30600000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.25200000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.17100000 0.24300000 ;
  END

END AO21x1_ASAP7_75t_L
MACRO TIELOx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN TIELOX1_ASAP7_75T_L 0 0 ;
 SIZE  0.16200000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.16200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.16200000 0.27900000 ;
    END
  END VDD

  PIN L
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09400000 0.02700000 0.14400000 0.04500000 ;
        RECT 0.12600000 0.04500000 0.14400000 0.18200000 ;
        RECT 0.06700000 0.18200000 0.14400000 0.20000000 ;
    END
  END L

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.09700000 0.09500000 0.11500000 ;
      RECT 0.01800000 0.11500000 0.03600000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.06800000 0.24300000 ;
  END

END TIELOx1_ASAP7_75t_L
MACRO DFFLQx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFLQX4_ASAP7_75T_L 0 0 ;
 SIZE  1.3500000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.35000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.35000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.12500000 0.06300000 1.25100000 0.08100000 ;
        RECT 1.20600000 0.08100000 1.22400000 0.18900000 ;
        RECT 1.12500000 0.18900000 1.25100000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.08300000 ;
      RECT 0.63900000 0.02700000 0.73800000 0.04500000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.08300000 ;
      RECT 0.66600000 0.10500000 0.68400000 0.14400000 ;
      RECT 0.93400000 0.06300000 0.98100000 0.08100000 ;
      RECT 0.96300000 0.08100000 0.98100000 0.10700000 ;
      RECT 0.96300000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.16400000 ;
      RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.06300000 ;
      RECT 0.18000000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
      RECT 1.01700000 0.06300000 1.06200000 0.08100000 ;
      RECT 1.04400000 0.08100000 1.06200000 0.10700000 ;
      RECT 1.04400000 0.10700000 1.11600000 0.12500000 ;
      RECT 1.09800000 0.12500000 1.11600000 0.14400000 ;
      RECT 1.04400000 0.12500000 1.06200000 0.18900000 ;
      RECT 1.01700000 0.18900000 1.06200000 0.20700000 ;
      RECT 0.54800000 0.06300000 0.58500000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.20900000 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.09000000 0.20700000 ;
      RECT 0.28800000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.07200000 0.20700000 0.09000000 0.22500000 ;
      RECT 0.28800000 0.20700000 0.30600000 0.22500000 ;
      RECT 0.07200000 0.22500000 0.30600000 0.24300000 ;
      RECT 0.39600000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.39600000 0.20700000 0.41400000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.41400000 0.24300000 ;
      RECT 0.50400000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.50400000 0.22500000 0.54100000 0.24300000 ;
      RECT 0.59200000 0.22500000 0.65700000 0.24300000 ;
      RECT 0.81900000 0.06300000 0.85600000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
      RECT 0.77400000 0.02700000 0.90000000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.45000000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.72000000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.58100000 0.20700000 ;
      RECT 0.51400000 0.22500000 0.62000000 0.24300000 ;
     LAYER V1 ;
      RECT 0.45000000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.55800000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.72000000 0.06300000 0.73800000 0.08100000 ;
      RECT 0.82800000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.93600000 0.06300000 0.95400000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.36000000 0.16200000 ;
      RECT 0.45000000 0.14400000 0.46800000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.46600000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.52100000 0.22500000 0.53900000 0.24300000 ;
      RECT 0.59400000 0.22500000 0.61200000 0.24300000 ;
  END

END DFFLQx4_ASAP7_75t_L
MACRO OR2x4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR2X4_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.02700000 0.25200000 0.04500000 ;
        RECT 0.23400000 0.04500000 0.25200000 0.06300000 ;
        RECT 0.23400000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.23400000 0.18900000 0.33300000 0.20700000 ;
        RECT 0.23400000 0.20700000 0.25200000 0.22500000 ;
        RECT 0.20700000 0.22500000 0.25200000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
  END

END OR2x4_ASAP7_75t_L
MACRO DECAPx4_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DECAPX4_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  OBS
     LAYER M1 ;
      RECT 0.23400000 0.06300000 0.49500000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.30600000 0.20700000 ;
  END

END DECAPx4_ASAP7_75t_L
MACRO AOI22xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI22XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END AOI22xp5_ASAP7_75t_L
MACRO AO21x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO21X2_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.30600000 0.04500000 ;
        RECT 0.28800000 0.04500000 0.30600000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.30600000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.06300000 0.25200000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.25200000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.17100000 0.24300000 ;
  END

END AO21x2_ASAP7_75t_L
MACRO INVx13_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX13_ASAP7_75T_L 0 0 ;
 SIZE  0.81 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.81000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.81000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.42300000 0.06300000 0.76500000 0.08100000 ;
        RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
        RECT 0.69300000 0.08100000 0.71100000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.76500000 0.20700000 ;
    END
  END Y

  OBS

  END

END INVx13_ASAP7_75t_L
MACRO AO221x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO221X2_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B2

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.47700000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
        RECT 0.47700000 0.18900000 0.52200000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.38700000 0.08100000 ;
      RECT 0.36900000 0.08100000 0.38700000 0.10700000 ;
      RECT 0.36900000 0.10700000 0.46800000 0.12500000 ;
      RECT 0.45000000 0.12500000 0.46800000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.11700000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.17100000 0.24300000 ;
      RECT 0.20700000 0.22500000 0.33300000 0.24300000 ;
  END

END AO221x2_ASAP7_75t_L
MACRO NOR4xp25_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR4XP25_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.04500000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A

  OBS

  END

END NOR4xp25_ASAP7_75t_L
MACRO ICGx5p33DC_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX5P33DC_ASAP7_75T_L 0 0 ;
 SIZE  2.5920000000000005 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 2.59200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 2.59200000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.09800000 0.12600000 1.11600000 0.16300000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.15200000 0.12600000 1.17000000 0.16300000 ;
    END
  END SE

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.61200000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.22500000 ;
        RECT 0.07200000 0.22500000 1.25100000 0.24300000 ;
        RECT 1.93500000 0.06300000 1.98000000 0.08100000 ;
        RECT 2.47500000 0.06300000 2.52000000 0.08100000 ;
        RECT 1.96200000 0.08100000 1.98000000 0.22500000 ;
        RECT 2.50200000 0.08100000 2.52000000 0.22500000 ;
        RECT 1.55500000 0.22500000 2.52000000 0.24300000 ;
       LAYER M2 ;
        RECT 1.23100000 0.22500000 1.57500000 0.24300000 ;
       LAYER V1 ;
        RECT 1.23100000 0.22500000 1.24900000 0.24300000 ;
        RECT 1.55700000 0.22500000 1.57500000 0.24300000 ;
    END
  END GCLK

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10500000 0.30600000 0.14400000 ;
        RECT 0.82800000 0.10500000 0.84600000 0.14400000 ;
        RECT 0.93600000 0.10500000 0.95400000 0.14400000 ;
        RECT 1.26000000 0.06300000 1.38600000 0.08100000 ;
        RECT 1.26000000 0.08100000 1.27800000 0.14400000 ;
        RECT 1.36800000 0.08100000 1.38600000 0.16400000 ;
        RECT 1.63800000 0.12600000 1.65600000 0.16400000 ;
        RECT 1.80000000 0.12600000 1.81800000 0.16400000 ;
        RECT 2.28600000 0.12600000 2.30400000 0.16400000 ;
       LAYER M2 ;
        RECT 0.28800000 0.10700000 1.27800000 0.12500000 ;
        RECT 1.36800000 0.14400000 2.30400000 0.16200000 ;
       LAYER V1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.82800000 0.10700000 0.84600000 0.12500000 ;
        RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
        RECT 1.26000000 0.10700000 1.27800000 0.12500000 ;
        RECT 1.36800000 0.14400000 1.38600000 0.16200000 ;
        RECT 1.63800000 0.14400000 1.65600000 0.16200000 ;
        RECT 1.80000000 0.14400000 1.81800000 0.16200000 ;
        RECT 2.28600000 0.14400000 2.30400000 0.16200000 ;
    END
  END CLK

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 1.69200000 0.06100000 1.71000000 0.14400000 ;
      RECT 2.04300000 0.06300000 2.16900000 0.08100000 ;
      RECT 2.12400000 0.08100000 2.14200000 0.14400000 ;
      RECT 1.85400000 0.02700000 2.41200000 0.04500000 ;
      RECT 1.85400000 0.04500000 1.87200000 0.06300000 ;
      RECT 1.80000000 0.06300000 1.87200000 0.08100000 ;
      RECT 1.85400000 0.08100000 1.87200000 0.14400000 ;
      RECT 2.23200000 0.04500000 2.25000000 0.14400000 ;
      RECT 2.39400000 0.04500000 2.41200000 0.14400000 ;
      RECT 1.52100000 0.06300000 1.55800000 0.08100000 ;
      RECT 1.53000000 0.08100000 1.54800000 0.16300000 ;
      RECT 0.23400000 0.06300000 0.27900000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.54900000 0.20700000 ;
      RECT 0.77400000 0.06300000 0.81900000 0.08100000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.18900000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.66600000 0.18900000 0.87300000 0.20700000 ;
      RECT 0.96300000 0.06300000 1.00800000 0.08100000 ;
      RECT 0.99000000 0.08100000 1.00800000 0.18900000 ;
      RECT 0.95700000 0.18900000 1.00800000 0.20700000 ;
      RECT 1.04400000 0.06300000 1.22400000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
      RECT 1.04400000 0.18900000 1.08900000 0.20700000 ;
      RECT 1.31400000 0.12600000 1.33200000 0.18900000 ;
      RECT 1.12300000 0.18900000 1.38600000 0.20700000 ;
      RECT 1.58400000 0.02700000 1.62900000 0.04500000 ;
      RECT 1.58400000 0.04500000 1.60200000 0.18900000 ;
      RECT 1.55500000 0.18900000 1.62900000 0.20700000 ;
      RECT 1.74600000 0.02700000 1.79100000 0.04500000 ;
      RECT 1.74600000 0.04500000 1.76400000 0.18900000 ;
      RECT 1.90800000 0.12600000 1.92600000 0.18900000 ;
      RECT 1.71900000 0.18900000 1.92600000 0.20700000 ;
      RECT 2.07000000 0.12600000 2.08800000 0.18900000 ;
      RECT 2.04300000 0.18900000 2.16900000 0.20700000 ;
      RECT 2.31300000 0.06300000 2.35800000 0.08100000 ;
      RECT 2.34000000 0.08100000 2.35800000 0.18900000 ;
      RECT 2.44800000 0.12600000 2.46600000 0.18900000 ;
      RECT 2.25900000 0.18900000 2.46600000 0.20700000 ;
      RECT 0.18000000 0.02700000 1.44000000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.14400000 ;
      RECT 0.34200000 0.04500000 0.36000000 0.14400000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.14400000 ;
      RECT 1.42200000 0.04500000 1.44000000 0.22500000 ;
      RECT 1.28700000 0.22500000 1.44000000 0.24300000 ;
      RECT 1.47600000 0.02700000 1.53500000 0.04500000 ;
      RECT 1.47600000 0.04500000 1.49400000 0.22500000 ;
      RECT 1.47600000 0.22500000 1.52100000 0.24300000 ;
     LAYER M2 ;
      RECT 1.53000000 0.06300000 1.82000000 0.08100000 ;
      RECT 0.96300000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.57500000 0.20700000 ;
     LAYER V1 ;
      RECT 1.53000000 0.06300000 1.54800000 0.08100000 ;
      RECT 1.69200000 0.06300000 1.71000000 0.08100000 ;
      RECT 1.80200000 0.06300000 1.82000000 0.08100000 ;
      RECT 0.96300000 0.18900000 0.98100000 0.20700000 ;
      RECT 1.12500000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.38400000 0.20700000 ;
      RECT 1.55700000 0.18900000 1.57500000 0.20700000 ;
  END

END ICGx5p33DC_ASAP7_75t_L
MACRO O2A1O1Ixp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN O2A1O1IXP33_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.30600000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.17100000 0.04500000 ;
      RECT 0.04500000 0.18900000 0.22500000 0.20700000 ;
  END

END O2A1O1Ixp33_ASAP7_75t_L
MACRO CKINVDCx9p33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX9P33_ASAP7_75T_L 0 0 ;
 SIZE  1.512 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.51200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.51200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.38700000 0.04500000 ;
        RECT 0.15300000 0.04500000 0.17100000 0.10700000 ;
        RECT 0.36900000 0.04500000 0.38700000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.17100000 0.12500000 ;
        RECT 0.36900000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.85500000 0.02700000 1.27800000 0.04500000 ;
        RECT 1.26000000 0.04500000 1.27800000 0.06300000 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
        RECT 1.26000000 0.06300000 1.41300000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.93600000 0.04500000 0.95400000 0.18900000 ;
        RECT 1.31400000 0.08100000 1.33200000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.14400000 0.20700000 ;
        RECT 0.80100000 0.18900000 0.98100000 0.20700000 ;
        RECT 1.28700000 0.18900000 1.41300000 0.20700000 ;
        RECT 0.12600000 0.20700000 0.14400000 0.22500000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.22500000 ;
        RECT 0.80100000 0.20700000 0.81900000 0.22500000 ;
        RECT 0.12600000 0.22500000 0.81900000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.14400000 ;
      RECT 0.63900000 0.06300000 0.76500000 0.08100000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.14400000 ;
      RECT 0.58500000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.58500000 0.04500000 0.60300000 0.10700000 ;
      RECT 0.80100000 0.04500000 0.81900000 0.10700000 ;
      RECT 0.55800000 0.10700000 0.60300000 0.12500000 ;
      RECT 0.80100000 0.10700000 0.84600000 0.12500000 ;
      RECT 0.55800000 0.12500000 0.57600000 0.14400000 ;
      RECT 0.82800000 0.12500000 0.84600000 0.14400000 ;
      RECT 1.07100000 0.06300000 1.19700000 0.08100000 ;
      RECT 1.15200000 0.08100000 1.17000000 0.14400000 ;
      RECT 0.28800000 0.12600000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.63900000 0.18900000 0.76500000 0.20700000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.18900000 ;
      RECT 1.07100000 0.18900000 1.19700000 0.20700000 ;
      RECT 0.99000000 0.12600000 1.00800000 0.14500000 ;
      RECT 1.26000000 0.12600000 1.27800000 0.14500000 ;
      RECT 0.99000000 0.14500000 1.03500000 0.16300000 ;
      RECT 1.23300000 0.14500000 1.27800000 0.16300000 ;
      RECT 1.01700000 0.16300000 1.03500000 0.22500000 ;
      RECT 1.23300000 0.16300000 1.25100000 0.22500000 ;
      RECT 1.01700000 0.22500000 1.25100000 0.24300000 ;
  END

END CKINVDCx9p33_ASAP7_75t_L
MACRO AO211x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO211X2_ASAP7_75T_L 0 0 ;
 SIZE  0.864 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.86400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.86400000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.12600000 0.33300000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.10700000 0.57600000 0.14400000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.74700000 0.06300000 0.79200000 0.08100000 ;
        RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
        RECT 0.74700000 0.18900000 0.79200000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.09900000 0.06300000 0.52200000 0.08100000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.14500000 ;
      RECT 0.61200000 0.14500000 0.73800000 0.16300000 ;
      RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
      RECT 0.61200000 0.16300000 0.63000000 0.18900000 ;
      RECT 0.50400000 0.18900000 0.63000000 0.20700000 ;
      RECT 0.31500000 0.22500000 0.60300000 0.24300000 ;
  END

END AO211x2_ASAP7_75t_L
MACRO XOR2x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XOR2X2_ASAP7_75T_L 0 0 ;
 SIZE  0.5940000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.38700000 0.04500000 ;
        RECT 0.26100000 0.04500000 0.27900000 0.06300000 ;
        RECT 0.12600000 0.06300000 0.27900000 0.08100000 ;
        RECT 0.36900000 0.04500000 0.38700000 0.10700000 ;
        RECT 0.36900000 0.10700000 0.41400000 0.12500000 ;
        RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
        RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.47700000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.22500000 ;
        RECT 0.47700000 0.22500000 0.52200000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.22500000 0.04500000 ;
      RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
      RECT 0.31500000 0.07600000 0.33300000 0.18900000 ;
      RECT 0.07200000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.01800000 0.06300000 0.06300000 0.08100000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.44100000 0.24300000 ;
  END

END XOR2x2_ASAP7_75t_L
MACRO DFFLQNx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFLQNX3_ASAP7_75T_L 0 0 ;
 SIZE  1.1880000000000004 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.18800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.18800000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.01700000 0.06300000 1.14300000 0.08100000 ;
        RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
        RECT 1.01700000 0.18900000 1.14300000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.42300000 0.02700000 0.46800000 0.04500000 ;
      RECT 0.45000000 0.04500000 0.46800000 0.08300000 ;
      RECT 0.66600000 0.10500000 0.68400000 0.14400000 ;
      RECT 0.93400000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.16400000 ;
      RECT 0.77400000 0.12600000 0.79200000 0.16400000 ;
      RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.06300000 ;
      RECT 0.18000000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.72000000 0.12600000 0.73800000 0.18900000 ;
      RECT 0.61200000 0.18900000 0.73800000 0.20700000 ;
      RECT 0.54800000 0.06300000 0.58500000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.20900000 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.11700000 0.20700000 ;
      RECT 0.26100000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.09900000 0.20700000 0.11700000 0.22500000 ;
      RECT 0.26100000 0.20700000 0.27900000 0.22500000 ;
      RECT 0.09900000 0.22500000 0.27900000 0.24300000 ;
      RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.42300000 0.20700000 0.44100000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.44100000 0.24300000 ;
      RECT 0.50400000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.50400000 0.22500000 0.54200000 0.24300000 ;
      RECT 0.59100000 0.22500000 0.65700000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.79200000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.06300000 ;
      RECT 0.77400000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.77400000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.77400000 0.20700000 0.79200000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.79200000 0.24300000 ;
      RECT 0.85500000 0.02700000 0.90000000 0.04500000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.45000000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.82800000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.77400000 0.14400000 0.90000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.58100000 0.20700000 ;
      RECT 0.51600000 0.22500000 0.61600000 0.24300000 ;
     LAYER V1 ;
      RECT 0.45000000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.55800000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.39600000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.82800000 0.10700000 0.84600000 0.12500000 ;
      RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.34200000 0.14400000 0.36000000 0.16200000 ;
      RECT 0.45000000 0.14400000 0.46800000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
      RECT 0.77400000 0.14400000 0.79200000 0.16200000 ;
      RECT 0.88200000 0.14400000 0.90000000 0.16200000 ;
      RECT 0.44800000 0.18900000 0.46600000 0.20700000 ;
      RECT 0.55800000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.52200000 0.22500000 0.54000000 0.24300000 ;
      RECT 0.59300000 0.22500000 0.61100000 0.24300000 ;
  END

END DFFLQNx3_ASAP7_75t_L
MACRO BUFx5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX5_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
        RECT 0.18000000 0.04500000 0.19800000 0.06300000 ;
        RECT 0.18000000 0.06300000 0.38700000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.38700000 0.20700000 ;
        RECT 0.20700000 0.20700000 0.22500000 0.22500000 ;
        RECT 0.15300000 0.22500000 0.22500000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx5_ASAP7_75t_L
MACRO AOI32xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI32XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.04500000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.26100000 0.18900000 0.36000000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.22500000 0.33300000 0.24300000 ;
  END

END AOI32xp33_ASAP7_75t_L
MACRO NOR3xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR3XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.17100000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END C

  OBS

  END

END NOR3xp33_ASAP7_75t_L
MACRO DHLx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DHLX3_ASAP7_75T_L 0 0 ;
 SIZE  0.9180000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.91800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.91800000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.69300000 0.06300000 0.81900000 0.08100000 ;
        RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
        RECT 0.69300000 0.18900000 0.81900000 0.20700000 ;
    END
  END Q

  OBS
     LAYER M1 ;
      RECT 0.66400000 0.10700000 0.73800000 0.12500000 ;
      RECT 0.72000000 0.12500000 0.73800000 0.14400000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.16400000 ;
      RECT 0.15300000 0.02700000 0.19800000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.06300000 ;
      RECT 0.18000000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.14400000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.15300000 0.18900000 0.19800000 0.20700000 ;
      RECT 0.01800000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.45000000 0.12600000 0.46800000 0.18900000 ;
      RECT 0.31500000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.22500000 ;
      RECT 0.31500000 0.20700000 0.33300000 0.22500000 ;
      RECT 0.01800000 0.22500000 0.33300000 0.24300000 ;
      RECT 0.42300000 0.02700000 0.52200000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.06300000 ;
      RECT 0.50400000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.50400000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.50400000 0.20700000 0.52200000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.52200000 0.24300000 ;
      RECT 0.58500000 0.02700000 0.63000000 0.04500000 ;
      RECT 0.61200000 0.04500000 0.63000000 0.22500000 ;
      RECT 0.58500000 0.22500000 0.63000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.55800000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.63000000 0.16200000 ;
     LAYER V1 ;
      RECT 0.55800000 0.10700000 0.57600000 0.12500000 ;
      RECT 0.66600000 0.10700000 0.68400000 0.12500000 ;
      RECT 0.50400000 0.14400000 0.52200000 0.16200000 ;
      RECT 0.61200000 0.14400000 0.63000000 0.16200000 ;
  END

END DHLx3_ASAP7_75t_L
MACRO OAI322xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI322XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.36900000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.15300000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END A3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.14400000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.04500000 0.06300000 0.27900000 0.08100000 ;
  END

END OAI322xp33_ASAP7_75t_L
MACRO AOI222xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI222XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.38700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END C1

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END C2

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END AOI222xp33_ASAP7_75t_L
MACRO DECAPx10_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DECAPX10_ASAP7_75T_L 0 0 ;
 SIZE  1.188 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.18800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.18800000 0.27900000 ;
    END
  END VDD

  OBS
     LAYER M1 ;
      RECT 0.55800000 0.06300000 1.14300000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.14400000 ;
      RECT 0.61200000 0.12600000 0.63000000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.63000000 0.20700000 ;
  END

END DECAPx10_ASAP7_75t_L
MACRO AND2x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND2X2_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.02700000 0.25200000 0.04500000 ;
        RECT 0.23400000 0.04500000 0.25200000 0.22500000 ;
        RECT 0.20700000 0.22500000 0.25200000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.19800000 0.20700000 ;
  END

END AND2x2_ASAP7_75t_L
MACRO NAND3x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND3X1_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.06300000 0.54900000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.44100000 0.20700000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.09900000 0.06300000 0.33300000 0.08100000 ;
  END

END NAND3x1_ASAP7_75t_L
MACRO AO22x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO22X2_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.42300000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.06300000 0.30600000 0.08100000 ;
      RECT 0.28800000 0.08100000 0.30600000 0.10700000 ;
      RECT 0.28800000 0.10700000 0.41400000 0.12500000 ;
      RECT 0.39600000 0.12500000 0.41400000 0.14400000 ;
      RECT 0.28800000 0.12500000 0.30600000 0.18900000 ;
      RECT 0.20700000 0.18900000 0.30600000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END AO22x2_ASAP7_75t_L
MACRO ICGx8DC_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX8DC_ASAP7_75T_L 0 0 ;
 SIZE  2.5920000000000005 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 2.59200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 2.59200000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.09800000 0.12600000 1.11600000 0.16300000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.15200000 0.12600000 1.17000000 0.16300000 ;
    END
  END SE

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.61200000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.22500000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.22500000 ;
        RECT 0.07200000 0.22500000 1.25100000 0.24300000 ;
        RECT 1.93500000 0.06300000 1.98000000 0.08100000 ;
        RECT 2.47500000 0.06300000 2.52000000 0.08100000 ;
        RECT 1.96200000 0.08100000 1.98000000 0.22500000 ;
        RECT 2.50200000 0.08100000 2.52000000 0.22500000 ;
        RECT 1.55500000 0.22500000 2.52000000 0.24300000 ;
       LAYER M2 ;
        RECT 1.23100000 0.22500000 1.57500000 0.24300000 ;
       LAYER V1 ;
        RECT 1.23100000 0.22500000 1.24900000 0.24300000 ;
        RECT 1.55700000 0.22500000 1.57500000 0.24300000 ;
    END
  END GCLK

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10500000 0.30600000 0.14400000 ;
        RECT 0.82800000 0.10500000 0.84600000 0.14400000 ;
        RECT 0.93600000 0.10500000 0.95400000 0.14400000 ;
        RECT 1.26000000 0.06300000 1.38600000 0.08100000 ;
        RECT 1.26000000 0.08100000 1.27800000 0.14400000 ;
        RECT 1.36800000 0.08100000 1.38600000 0.16400000 ;
       LAYER M2 ;
        RECT 0.28800000 0.10700000 1.27800000 0.12500000 ;
       LAYER V1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.82800000 0.10700000 0.84600000 0.12500000 ;
        RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
        RECT 1.26000000 0.10700000 1.27800000 0.12500000 ;
    END
  END CLK

  OBS
     LAYER M1 ;
      RECT 1.52100000 0.06300000 1.55800000 0.08100000 ;
      RECT 1.53000000 0.08100000 1.54800000 0.12500000 ;
      RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 2.04300000 0.06300000 2.16900000 0.08100000 ;
      RECT 2.12400000 0.08100000 2.14200000 0.14400000 ;
      RECT 1.69200000 0.02700000 2.41200000 0.04500000 ;
      RECT 1.69200000 0.04500000 1.71000000 0.06300000 ;
      RECT 1.63800000 0.06300000 1.71000000 0.08100000 ;
      RECT 1.69200000 0.08100000 1.71000000 0.14400000 ;
      RECT 1.85400000 0.04500000 1.87200000 0.14400000 ;
      RECT 2.23200000 0.04500000 2.25000000 0.14400000 ;
      RECT 2.39400000 0.04500000 2.41200000 0.14400000 ;
      RECT 1.63800000 0.12600000 1.65600000 0.16400000 ;
      RECT 1.80000000 0.12600000 1.81800000 0.16400000 ;
      RECT 2.28600000 0.12600000 2.30400000 0.16400000 ;
      RECT 0.23400000 0.06300000 0.27900000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.54900000 0.20700000 ;
      RECT 0.77400000 0.06300000 0.81900000 0.08100000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.18900000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.18900000 ;
      RECT 0.66600000 0.18900000 0.87300000 0.20700000 ;
      RECT 0.96300000 0.06300000 1.00800000 0.08100000 ;
      RECT 0.99000000 0.08100000 1.00800000 0.18900000 ;
      RECT 0.95500000 0.18900000 1.00800000 0.20700000 ;
      RECT 1.04400000 0.06300000 1.22400000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
      RECT 1.04400000 0.18900000 1.08900000 0.20700000 ;
      RECT 1.31400000 0.12600000 1.33200000 0.18900000 ;
      RECT 1.12300000 0.18900000 1.38600000 0.20700000 ;
      RECT 1.58400000 0.02700000 1.62900000 0.04500000 ;
      RECT 1.58400000 0.04500000 1.60200000 0.18900000 ;
      RECT 1.55500000 0.18900000 1.62900000 0.20700000 ;
      RECT 1.74600000 0.06300000 1.79100000 0.08100000 ;
      RECT 1.74600000 0.08100000 1.76400000 0.18900000 ;
      RECT 1.90800000 0.12600000 1.92600000 0.18900000 ;
      RECT 1.71900000 0.18900000 1.92600000 0.20700000 ;
      RECT 2.07000000 0.12600000 2.08800000 0.18900000 ;
      RECT 2.04300000 0.18900000 2.16900000 0.20700000 ;
      RECT 2.31300000 0.06300000 2.35800000 0.08100000 ;
      RECT 2.34000000 0.08100000 2.35800000 0.18900000 ;
      RECT 2.44800000 0.12600000 2.46600000 0.18900000 ;
      RECT 2.25900000 0.18900000 2.46600000 0.20700000 ;
      RECT 0.18000000 0.02700000 1.44000000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.14400000 ;
      RECT 0.34200000 0.04500000 0.36000000 0.14400000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.14400000 ;
      RECT 1.42200000 0.04500000 1.44000000 0.22500000 ;
      RECT 1.28700000 0.22500000 1.44000000 0.24300000 ;
      RECT 1.47600000 0.02700000 1.53900000 0.04500000 ;
      RECT 1.47600000 0.04500000 1.49400000 0.22500000 ;
      RECT 1.47600000 0.22500000 1.52100000 0.24300000 ;
     LAYER M2 ;
      RECT 1.53000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14400000 2.30400000 0.16200000 ;
      RECT 0.96300000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.57500000 0.20700000 ;
     LAYER V1 ;
      RECT 1.53000000 0.06300000 1.54800000 0.08100000 ;
      RECT 1.64000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14400000 1.38600000 0.16200000 ;
      RECT 1.63800000 0.14400000 1.65600000 0.16200000 ;
      RECT 1.80000000 0.14400000 1.81800000 0.16200000 ;
      RECT 2.28600000 0.14400000 2.30400000 0.16200000 ;
      RECT 0.96300000 0.18900000 0.98100000 0.20700000 ;
      RECT 1.12500000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.38400000 0.20700000 ;
      RECT 1.55700000 0.18900000 1.57500000 0.20700000 ;
  END

END ICGx8DC_ASAP7_75t_L
MACRO NOR5xp2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR5XP2_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.33300000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END D

  PIN E
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END E

  OBS

  END

END NOR5xp2_ASAP7_75t_L
MACRO XOR2xp5_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XOR2XP5_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.14500000 ;
        RECT 0.28800000 0.12600000 0.30600000 0.14500000 ;
        RECT 0.12600000 0.14500000 0.30600000 0.16300000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.26100000 0.02700000 0.46800000 0.04500000 ;
        RECT 0.45000000 0.04500000 0.46800000 0.22500000 ;
        RECT 0.42300000 0.22500000 0.46800000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.02700000 0.11700000 0.04500000 ;
      RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.41400000 0.20700000 ;
      RECT 0.26100000 0.22500000 0.38700000 0.24300000 ;
  END

END XOR2xp5_ASAP7_75t_L
MACRO AO222x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO222X2_ASAP7_75T_L 0 0 ;
 SIZE  0.648 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.64800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.64800000 0.27900000 ;
    END
  END VDD

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END C1

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END C2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END A2

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.53100000 0.02700000 0.57600000 0.04500000 ;
        RECT 0.55800000 0.04500000 0.57600000 0.18900000 ;
        RECT 0.53100000 0.18900000 0.57600000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.52200000 0.08100000 ;
      RECT 0.50400000 0.08100000 0.52200000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.11700000 0.20700000 ;
      RECT 0.20700000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END AO222x2_ASAP7_75t_L
MACRO MAJx3_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN MAJX3_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.30600000 0.08100000 ;
        RECT 0.15300000 0.08100000 0.17100000 0.10700000 ;
        RECT 0.12600000 0.10700000 0.17100000 0.12500000 ;
        RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END C

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.36900000 0.06300000 0.49500000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.22500000 ;
        RECT 0.36900000 0.22500000 0.49500000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.34200000 0.12600000 0.36000000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.36000000 0.20700000 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END MAJx3_ASAP7_75t_L
MACRO OR5x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR5X2_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END D

  PIN E
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END E

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.36900000 0.02700000 0.41400000 0.04500000 ;
        RECT 0.39600000 0.04500000 0.41400000 0.18900000 ;
        RECT 0.36900000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.36000000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
  END

END OR5x2_ASAP7_75t_L
MACRO AO32x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO32X1_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.02700000 0.06300000 0.04500000 ;
        RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  OBS
     LAYER M1 ;
      RECT 0.07200000 0.06300000 0.41400000 0.08100000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
      RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
      RECT 0.31500000 0.18900000 0.41400000 0.20700000 ;
      RECT 0.15300000 0.22500000 0.38700000 0.24300000 ;
  END

END AO32x1_ASAP7_75t_L
MACRO AOI22x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI22X1_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.04500000 0.02700000 0.46800000 0.04500000 ;
        RECT 0.45000000 0.04500000 0.46800000 0.06300000 ;
        RECT 0.45000000 0.06300000 0.52200000 0.08100000 ;
        RECT 0.50400000 0.08100000 0.52200000 0.18900000 ;
        RECT 0.31500000 0.18900000 0.52200000 0.20700000 ;
    END
  END Y

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.14500000 ;
        RECT 0.20700000 0.14500000 0.25200000 0.16300000 ;
        RECT 0.07200000 0.12600000 0.09000000 0.18900000 ;
        RECT 0.20700000 0.16300000 0.22500000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.22500000 0.20700000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.10700000 0.17100000 0.14400000 ;
    END
  END B1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.06300000 0.41400000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.10700000 ;
        RECT 0.39600000 0.10700000 0.46800000 0.12500000 ;
        RECT 0.28800000 0.08100000 0.30600000 0.14400000 ;
        RECT 0.45000000 0.12500000 0.46800000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.22500000 0.49500000 0.24300000 ;
  END

END AOI22x1_ASAP7_75t_L
MACRO BUFx10_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX10_ASAP7_75T_L 0 0 ;
 SIZE  0.756 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.75600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.75600000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.65700000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14500000 ;
      RECT 0.18000000 0.12600000 0.19800000 0.14500000 ;
      RECT 0.12600000 0.14500000 0.19800000 0.16300000 ;
      RECT 0.12600000 0.16300000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx10_ASAP7_75t_L
MACRO ICGx4DC_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN ICGX4DC_ASAP7_75T_L 0 0 ;
 SIZE  2.5920000000000005 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 2.59200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 2.59200000 0.27900000 ;
    END
  END VDD

  PIN ENA
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.09800000 0.12600000 1.11600000 0.16300000 ;
    END
  END ENA

  PIN SE
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.15200000 0.12600000 1.17000000 0.16300000 ;
    END
  END SE

  PIN GCLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.61200000 0.06300000 0.65700000 0.08100000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.22500000 ;
        RECT 0.61200000 0.08100000 0.63000000 0.22500000 ;
        RECT 0.07200000 0.22500000 1.25100000 0.24300000 ;
        RECT 2.47500000 0.02700000 2.52000000 0.04500000 ;
        RECT 1.93500000 0.06300000 1.98000000 0.08100000 ;
        RECT 1.96200000 0.08100000 1.98000000 0.22500000 ;
        RECT 2.50200000 0.04500000 2.52000000 0.22500000 ;
        RECT 1.57800000 0.22500000 2.52000000 0.24300000 ;
       LAYER M2 ;
        RECT 1.23100000 0.22500000 1.59900000 0.24300000 ;
       LAYER V1 ;
        RECT 1.23100000 0.22500000 1.24900000 0.24300000 ;
        RECT 1.58100000 0.22500000 1.59900000 0.24300000 ;
    END
  END GCLK

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10500000 0.30600000 0.14400000 ;
        RECT 0.77400000 0.10500000 0.79200000 0.14400000 ;
        RECT 0.93600000 0.10500000 0.95400000 0.14400000 ;
        RECT 1.26000000 0.06300000 1.38600000 0.08100000 ;
        RECT 1.26000000 0.08100000 1.27800000 0.14400000 ;
        RECT 1.36800000 0.08100000 1.38600000 0.16400000 ;
       LAYER M2 ;
        RECT 0.28800000 0.10700000 1.27800000 0.12500000 ;
       LAYER V1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.12500000 ;
        RECT 0.77400000 0.10700000 0.79200000 0.12500000 ;
        RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
        RECT 1.26000000 0.10700000 1.27800000 0.12500000 ;
    END
  END CLK

  OBS
     LAYER M1 ;
      RECT 1.52100000 0.06300000 1.55800000 0.08100000 ;
      RECT 1.53000000 0.08100000 1.54800000 0.12500000 ;
      RECT 0.42300000 0.06300000 0.54900000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 2.04300000 0.06300000 2.16900000 0.08100000 ;
      RECT 2.12400000 0.08100000 2.14200000 0.14400000 ;
      RECT 1.71900000 0.02700000 2.41200000 0.04500000 ;
      RECT 1.71900000 0.04500000 1.73700000 0.06300000 ;
      RECT 1.63800000 0.06300000 1.73700000 0.08100000 ;
      RECT 1.69200000 0.08100000 1.71000000 0.14400000 ;
      RECT 1.85400000 0.04500000 1.87200000 0.14400000 ;
      RECT 2.23200000 0.04500000 2.25000000 0.14400000 ;
      RECT 2.39400000 0.04500000 2.41200000 0.14400000 ;
      RECT 1.63800000 0.12600000 1.65600000 0.16400000 ;
      RECT 1.74600000 0.12600000 1.76400000 0.16400000 ;
      RECT 2.28600000 0.12600000 2.30400000 0.16400000 ;
      RECT 0.23400000 0.06300000 0.27900000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.18900000 ;
      RECT 0.12600000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.50400000 0.12600000 0.52200000 0.18900000 ;
      RECT 0.42300000 0.18900000 0.54900000 0.20700000 ;
      RECT 0.80100000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.18900000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.66600000 0.18900000 0.87300000 0.20700000 ;
      RECT 0.96300000 0.06300000 1.00800000 0.08100000 ;
      RECT 0.99000000 0.08100000 1.00800000 0.18900000 ;
      RECT 0.95700000 0.18900000 1.00800000 0.20700000 ;
      RECT 1.04400000 0.06300000 1.22400000 0.08100000 ;
      RECT 1.20600000 0.08100000 1.22400000 0.14400000 ;
      RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
      RECT 1.04400000 0.18900000 1.08900000 0.20700000 ;
      RECT 1.31400000 0.12600000 1.33200000 0.18900000 ;
      RECT 1.12300000 0.18900000 1.38600000 0.20700000 ;
      RECT 1.58400000 0.02700000 1.62900000 0.04500000 ;
      RECT 1.58400000 0.04500000 1.60200000 0.18900000 ;
      RECT 1.53000000 0.18900000 1.62900000 0.20700000 ;
      RECT 1.77300000 0.06300000 1.81800000 0.08100000 ;
      RECT 1.80000000 0.08100000 1.81800000 0.18900000 ;
      RECT 1.90800000 0.12600000 1.92600000 0.18900000 ;
      RECT 1.71900000 0.18900000 1.92600000 0.20700000 ;
      RECT 2.07000000 0.12600000 2.08800000 0.18900000 ;
      RECT 2.04300000 0.18900000 2.16900000 0.20700000 ;
      RECT 2.31300000 0.06300000 2.35800000 0.08100000 ;
      RECT 2.34000000 0.08100000 2.35800000 0.18900000 ;
      RECT 2.44800000 0.12600000 2.46600000 0.18900000 ;
      RECT 2.25900000 0.18900000 2.46600000 0.20700000 ;
      RECT 0.18000000 0.02700000 1.44000000 0.04500000 ;
      RECT 0.18000000 0.04500000 0.19800000 0.14400000 ;
      RECT 0.34200000 0.04500000 0.36000000 0.14400000 ;
      RECT 0.72000000 0.04500000 0.73800000 0.14400000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.14400000 ;
      RECT 1.42200000 0.04500000 1.44000000 0.22500000 ;
      RECT 1.28700000 0.22500000 1.44000000 0.24300000 ;
      RECT 1.47600000 0.02700000 1.54300000 0.04500000 ;
      RECT 1.47600000 0.04500000 1.49400000 0.22500000 ;
      RECT 1.47600000 0.22500000 1.52100000 0.24300000 ;
     LAYER M2 ;
      RECT 1.53000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14400000 2.30400000 0.16200000 ;
      RECT 0.96300000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.55000000 0.20700000 ;
     LAYER V1 ;
      RECT 1.53000000 0.06300000 1.54800000 0.08100000 ;
      RECT 1.64000000 0.06300000 1.65800000 0.08100000 ;
      RECT 1.36800000 0.14400000 1.38600000 0.16200000 ;
      RECT 1.63800000 0.14400000 1.65600000 0.16200000 ;
      RECT 1.74600000 0.14400000 1.76400000 0.16200000 ;
      RECT 2.28600000 0.14400000 2.30400000 0.16200000 ;
      RECT 0.96300000 0.18900000 0.98100000 0.20700000 ;
      RECT 1.12500000 0.18900000 1.14300000 0.20700000 ;
      RECT 1.36600000 0.18900000 1.38400000 0.20700000 ;
      RECT 1.53200000 0.18900000 1.55000000 0.20700000 ;
  END

END ICGx4DC_ASAP7_75t_L
MACRO AO333x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO333X2_ASAP7_75T_L 0 0 ;
 SIZE  0.7020000000000001 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.70200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.70200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.02700000 0.11700000 0.04500000 ;
        RECT 0.07200000 0.04500000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END B1

  PIN C3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END C3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.12600000 0.57600000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.12600000 0.63000000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.20700000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.12600000 0.06300000 0.68400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14400000 ;
      RECT 0.66600000 0.08100000 0.68400000 0.18900000 ;
      RECT 0.53100000 0.18900000 0.68400000 0.20700000 ;
      RECT 0.36900000 0.22500000 0.60300000 0.24300000 ;
  END

END AO333x2_ASAP7_75t_L
MACRO OAI21xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI21XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.27 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.27000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.27000000 0.27900000 ;
    END
  END VDD

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.17100000 0.20700000 ;
    END
  END Y

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.02700000 0.17100000 0.04500000 ;
  END

END OAI21xp33_ASAP7_75t_L
MACRO NOR2xp67_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR2XP67_ASAP7_75T_L 0 0 ;
 SIZE  0.32400000000000007 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.06300000 0.17100000 0.18900000 ;
        RECT 0.15300000 0.18900000 0.22500000 0.20700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.12600000 0.11700000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.12600000 0.22500000 0.16300000 ;
    END
  END B

  OBS
     LAYER M1 ;
      RECT 0.04500000 0.22500000 0.27900000 0.24300000 ;
  END

END NOR2xp67_ASAP7_75t_L
MACRO NAND4xp75_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NAND4XP75_ASAP7_75T_L 0 0 ;
 SIZE  0.756 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.75600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.75600000 0.27900000 ;
    END
  END VDD

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.12600000 0.11700000 0.16300000 ;
    END
  END D

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.55800000 0.06300000 0.71100000 0.08100000 ;
        RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.65700000 0.20700000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.47700000 0.12600000 0.49500000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.63900000 0.12600000 0.65700000 0.16300000 ;
    END
  END A

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.33300000 0.04500000 ;
      RECT 0.42300000 0.02700000 0.65700000 0.04500000 ;
      RECT 0.26100000 0.06300000 0.49500000 0.08100000 ;
  END

END NAND4xp75_ASAP7_75t_L
MACRO AOI331xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI331XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.486 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.48600000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.48600000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.46800000 0.08100000 ;
        RECT 0.45000000 0.08100000 0.46800000 0.18900000 ;
        RECT 0.42300000 0.18900000 0.46800000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.26100000 0.22500000 0.38700000 0.24300000 ;
  END

END AOI331xp33_ASAP7_75t_L
MACRO OR2x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR2X2_ASAP7_75T_L 0 0 ;
 SIZE  0.324 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.32400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.32400000 0.27900000 ;
    END
  END VDD

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.02700000 0.25200000 0.04500000 ;
        RECT 0.23400000 0.04500000 0.25200000 0.22500000 ;
        RECT 0.20700000 0.22500000 0.25200000 0.24300000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.04500000 0.18900000 0.19800000 0.20700000 ;
  END

END OR2x2_ASAP7_75t_L
MACRO AO332x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AO332X1_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.01800000 0.02700000 0.06300000 0.04500000 ;
        RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
        RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
    END
  END Y

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END B3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.15300000 0.18900000 0.38700000 0.20700000 ;
      RECT 0.07200000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.47700000 0.18900000 0.57600000 0.20700000 ;
      RECT 0.31500000 0.22500000 0.54900000 0.24300000 ;
  END

END AO332x1_ASAP7_75t_L
MACRO AOI333xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI333XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.594 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN C3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END C3

  PIN C2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END C2

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.57600000 0.08100000 ;
        RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
        RECT 0.42300000 0.18900000 0.57600000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END B1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END B2

  PIN B3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16300000 ;
    END
  END B3

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.12600000 0.41400000 0.16300000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.12600000 0.46800000 0.16300000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END A1

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.18900000 0.33300000 0.20700000 ;
      RECT 0.26100000 0.22500000 0.49500000 0.24300000 ;
  END

END AOI333xp33_ASAP7_75t_L
MACRO OA22x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA22X2_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.34200000 0.10700000 0.36000000 0.14400000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.39600000 0.10700000 0.41400000 0.14400000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.45000000 0.10700000 0.46800000 0.14400000 ;
    END
  END B1

  OBS
     LAYER M1 ;
      RECT 0.26100000 0.02700000 0.49500000 0.04500000 ;
      RECT 0.23400000 0.06300000 0.33300000 0.08100000 ;
      RECT 0.23400000 0.08100000 0.25200000 0.10700000 ;
      RECT 0.12600000 0.10700000 0.25200000 0.12500000 ;
      RECT 0.12600000 0.12500000 0.14400000 0.14400000 ;
      RECT 0.23400000 0.12500000 0.25200000 0.18900000 ;
      RECT 0.23400000 0.18900000 0.38700000 0.20700000 ;
  END

END OA22x2_ASAP7_75t_L
MACRO INVxp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVXP33_ASAP7_75T_L 0 0 ;
 SIZE  0.162 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.16200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.16200000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.09900000 0.02700000 0.14400000 0.04500000 ;
        RECT 0.12600000 0.04500000 0.14400000 0.22500000 ;
        RECT 0.09900000 0.22500000 0.14400000 0.24300000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  OBS

  END

END INVxp33_ASAP7_75t_L
MACRO DFFLQNx1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN DFFLQNX1_ASAP7_75T_L 0 0 ;
 SIZE  1.0800000000000003 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 1.08000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 1.08000000 0.27900000 ;
    END
  END VDD

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END D

  PIN QN
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 1.01700000 0.06300000 1.06200000 0.08100000 ;
        RECT 1.04400000 0.08100000 1.06200000 0.18900000 ;
        RECT 1.01700000 0.18900000 1.06200000 0.20700000 ;
    END
  END QN

  OBS
     LAYER M1 ;
      RECT 0.39600000 0.02700000 0.45300000 0.04500000 ;
      RECT 0.39600000 0.04500000 0.41400000 0.06300000 ;
      RECT 0.39600000 0.06300000 0.45400000 0.08100000 ;
      RECT 0.45000000 0.10600000 0.46800000 0.14400000 ;
      RECT 0.61200000 0.06300000 0.73800000 0.08100000 ;
      RECT 0.61200000 0.08100000 0.63000000 0.14400000 ;
      RECT 0.72000000 0.08100000 0.73800000 0.14400000 ;
      RECT 0.93400000 0.10700000 1.00800000 0.12500000 ;
      RECT 0.99000000 0.12500000 1.00800000 0.14400000 ;
      RECT 0.77400000 0.12600000 0.79200000 0.16400000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.16500000 ;
      RECT 0.09900000 0.02700000 0.27900000 0.04500000 ;
      RECT 0.09900000 0.04500000 0.11700000 0.06300000 ;
      RECT 0.26100000 0.04500000 0.27900000 0.06300000 ;
      RECT 0.01800000 0.06300000 0.11700000 0.08100000 ;
      RECT 0.26100000 0.06300000 0.36000000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.14400000 0.20700000 ;
      RECT 0.54900000 0.06300000 0.58600000 0.08100000 ;
      RECT 0.55800000 0.08100000 0.57600000 0.18900000 ;
      RECT 0.55800000 0.18900000 0.60300000 0.20700000 ;
      RECT 0.15300000 0.06300000 0.19800000 0.08100000 ;
      RECT 0.18000000 0.08100000 0.19800000 0.18900000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.41400000 0.20700000 ;
      RECT 0.18000000 0.20700000 0.19800000 0.22500000 ;
      RECT 0.15300000 0.22500000 0.19800000 0.24300000 ;
      RECT 0.45000000 0.18700000 0.46800000 0.22500000 ;
      RECT 0.36900000 0.22500000 0.46800000 0.24300000 ;
      RECT 0.50400000 0.02700000 0.60300000 0.04500000 ;
      RECT 0.50400000 0.04500000 0.52200000 0.22500000 ;
      RECT 0.50400000 0.22500000 0.60300000 0.24300000 ;
      RECT 0.63900000 0.02700000 0.79200000 0.04500000 ;
      RECT 0.77400000 0.04500000 0.79200000 0.06300000 ;
      RECT 0.77400000 0.06300000 0.84600000 0.08100000 ;
      RECT 0.82800000 0.08100000 0.84600000 0.18900000 ;
      RECT 0.72000000 0.18900000 0.84600000 0.20700000 ;
      RECT 0.72000000 0.20700000 0.73800000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.73800000 0.24300000 ;
      RECT 0.85500000 0.02700000 0.90000000 0.04500000 ;
      RECT 0.88200000 0.04500000 0.90000000 0.22500000 ;
      RECT 0.85500000 0.22500000 0.90000000 0.24300000 ;
     LAYER M2 ;
      RECT 0.42100000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.82800000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.34200000 0.10800000 0.63000000 0.12600000 ;
      RECT 0.77400000 0.14400000 0.90000000 0.16200000 ;
      RECT 0.39600000 0.14500000 0.68400000 0.16300000 ;
      RECT 0.45000000 0.18900000 0.60100000 0.20700000 ;
     LAYER V1 ;
      RECT 0.42100000 0.06300000 0.43900000 0.08100000 ;
      RECT 0.55800000 0.06300000 0.57600000 0.08100000 ;
      RECT 0.82800000 0.10700000 0.84600000 0.12500000 ;
      RECT 0.93600000 0.10700000 0.95400000 0.12500000 ;
      RECT 0.34200000 0.10800000 0.36000000 0.12600000 ;
      RECT 0.45000000 0.10800000 0.46800000 0.12600000 ;
      RECT 0.61200000 0.10800000 0.63000000 0.12600000 ;
      RECT 0.77400000 0.14400000 0.79200000 0.16200000 ;
      RECT 0.88200000 0.14400000 0.90000000 0.16200000 ;
      RECT 0.39600000 0.14500000 0.41400000 0.16300000 ;
      RECT 0.66600000 0.14500000 0.68400000 0.16300000 ;
      RECT 0.45000000 0.18900000 0.46800000 0.20700000 ;
      RECT 0.58300000 0.18900000 0.60100000 0.20700000 ;
  END

END DFFLQNx1_ASAP7_75t_L
MACRO CKINVDCx20_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CKINVDCX20_ASAP7_75T_L 0 0 ;
 SIZE  2.052 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 2.05200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 2.05200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.14500000 ;
        RECT 0.50400000 0.12600000 0.52200000 0.14500000 ;
        RECT 0.23400000 0.14500000 0.27900000 0.16300000 ;
        RECT 0.47700000 0.14500000 0.52200000 0.16300000 ;
        RECT 0.26100000 0.16300000 0.27900000 0.22500000 ;
        RECT 0.47700000 0.16300000 0.49500000 0.22500000 ;
        RECT 0.26100000 0.22500000 0.49500000 0.24300000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.15300000 0.02700000 1.95300000 0.04500000 ;
        RECT 0.15300000 0.04500000 0.17100000 0.06300000 ;
        RECT 0.09900000 0.06300000 0.17100000 0.08100000 ;
        RECT 0.15300000 0.08100000 0.17100000 0.18900000 ;
        RECT 0.55800000 0.04500000 0.57600000 0.18900000 ;
        RECT 0.99000000 0.04500000 1.00800000 0.18900000 ;
        RECT 1.44900000 0.04500000 1.46700000 0.18900000 ;
        RECT 1.85400000 0.04500000 1.87200000 0.18900000 ;
        RECT 0.09900000 0.18900000 0.22500000 0.20700000 ;
        RECT 0.53100000 0.18900000 0.65700000 0.20700000 ;
        RECT 0.96300000 0.18900000 1.08900000 0.20700000 ;
        RECT 1.39500000 0.18900000 1.52100000 0.20700000 ;
        RECT 1.82700000 0.18900000 1.95300000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.31500000 0.06300000 0.44100000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.74700000 0.06300000 0.87300000 0.08100000 ;
      RECT 0.77400000 0.08100000 0.79200000 0.14400000 ;
      RECT 1.17900000 0.06300000 1.30500000 0.08100000 ;
      RECT 1.26000000 0.08100000 1.27800000 0.14400000 ;
      RECT 1.61100000 0.06300000 1.73700000 0.08100000 ;
      RECT 1.69200000 0.08100000 1.71000000 0.14400000 ;
      RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
      RECT 0.31500000 0.18900000 0.44100000 0.20700000 ;
      RECT 0.82800000 0.12600000 0.84600000 0.18900000 ;
      RECT 0.74700000 0.18900000 0.87300000 0.20700000 ;
      RECT 1.20600000 0.12600000 1.22400000 0.18900000 ;
      RECT 1.17900000 0.18900000 1.30500000 0.20700000 ;
      RECT 1.63800000 0.12600000 1.65600000 0.18900000 ;
      RECT 1.61100000 0.18900000 1.73700000 0.20700000 ;
      RECT 0.66600000 0.12600000 0.68400000 0.14500000 ;
      RECT 0.93600000 0.12600000 0.95400000 0.14500000 ;
      RECT 0.66600000 0.14500000 0.71100000 0.16300000 ;
      RECT 0.90900000 0.14500000 0.95400000 0.16300000 ;
      RECT 0.69300000 0.16300000 0.71100000 0.22500000 ;
      RECT 0.90900000 0.16300000 0.92700000 0.22500000 ;
      RECT 0.69300000 0.22500000 0.92700000 0.24300000 ;
      RECT 1.09800000 0.12600000 1.11600000 0.14500000 ;
      RECT 1.36800000 0.12600000 1.38600000 0.14500000 ;
      RECT 1.09800000 0.14500000 1.14300000 0.16300000 ;
      RECT 1.34100000 0.14500000 1.38600000 0.16300000 ;
      RECT 1.12500000 0.16300000 1.14300000 0.22500000 ;
      RECT 1.34100000 0.16300000 1.35900000 0.22500000 ;
      RECT 1.12500000 0.22500000 1.35900000 0.24300000 ;
      RECT 1.53000000 0.12600000 1.54800000 0.14500000 ;
      RECT 1.80000000 0.12600000 1.81800000 0.14500000 ;
      RECT 1.53000000 0.14500000 1.57500000 0.16300000 ;
      RECT 1.77300000 0.14500000 1.81800000 0.16300000 ;
      RECT 1.55700000 0.16300000 1.57500000 0.22500000 ;
      RECT 1.77300000 0.16300000 1.79100000 0.22500000 ;
      RECT 1.55700000 0.22500000 1.79100000 0.24300000 ;
  END

END CKINVDCx20_ASAP7_75t_L
MACRO OAI311xp33_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI311XP33_ASAP7_75T_L 0 0 ;
 SIZE  0.378 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.37800000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.37800000 0.27900000 ;
    END
  END VDD

  PIN A3
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A3

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.10700000 0.14400000 0.14400000 ;
    END
  END A2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.10700000 0.19800000 0.14400000 ;
    END
  END A1

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.06300000 0.36000000 0.08100000 ;
        RECT 0.34200000 0.08100000 0.36000000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.36000000 0.20700000 ;
    END
  END Y

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.10700000 0.25200000 0.14400000 ;
    END
  END B1

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.10700000 0.30600000 0.14400000 ;
    END
  END C1

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.02700000 0.22500000 0.04500000 ;
  END

END OAI311xp33_ASAP7_75t_L
MACRO OA221x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OA221X2_ASAP7_75T_L 0 0 ;
 SIZE  0.8640000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.86400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.86400000 0.27900000 ;
    END
  END VDD

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.06300000 0.11700000 0.08100000 ;
        RECT 0.07200000 0.08100000 0.09000000 0.18900000 ;
        RECT 0.07200000 0.18900000 0.11700000 0.20700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END A1

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.31500000 0.12600000 0.33300000 0.16300000 ;
    END
  END A2

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.50400000 0.12600000 0.52200000 0.16300000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.61200000 0.12600000 0.63000000 0.16300000 ;
    END
  END B1

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.77400000 0.10700000 0.79200000 0.14400000 ;
    END
  END C

  OBS
     LAYER M1 ;
      RECT 0.47700000 0.02700000 0.81900000 0.04500000 ;
      RECT 0.20700000 0.06300000 0.65700000 0.08100000 ;
      RECT 0.72000000 0.06300000 0.76500000 0.08100000 ;
      RECT 0.12600000 0.12600000 0.14400000 0.14500000 ;
      RECT 0.12600000 0.14500000 0.19800000 0.16300000 ;
      RECT 0.18000000 0.16300000 0.19800000 0.18900000 ;
      RECT 0.72000000 0.08100000 0.73800000 0.18900000 ;
      RECT 0.18000000 0.18900000 0.76500000 0.20700000 ;
  END

END OA221x2_ASAP7_75t_L
MACRO BUFx6f_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN BUFX6F_ASAP7_75T_L 0 0 ;
 SIZE  0.54 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.54000000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.54000000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.10700000 0.09000000 0.14400000 ;
    END
  END A

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.20700000 0.06300000 0.44100000 0.08100000 ;
        RECT 0.39600000 0.08100000 0.41400000 0.18900000 ;
        RECT 0.20700000 0.18900000 0.44100000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.09900000 0.06300000 0.14400000 0.08100000 ;
      RECT 0.12600000 0.08100000 0.14400000 0.14500000 ;
      RECT 0.18000000 0.12600000 0.19800000 0.14500000 ;
      RECT 0.12600000 0.14500000 0.19800000 0.16300000 ;
      RECT 0.12600000 0.16300000 0.14400000 0.18900000 ;
      RECT 0.09900000 0.18900000 0.14400000 0.20700000 ;
  END

END BUFx6f_ASAP7_75t_L
MACRO OR5x1_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OR5X1_ASAP7_75T_L 0 0 ;
 SIZE  0.432 BY 0.27 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.43200000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.43200000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.07200000 0.12600000 0.09000000 0.16300000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.16300000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.16300000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.23400000 0.12600000 0.25200000 0.16300000 ;
    END
  END D

  PIN E
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.28800000 0.12600000 0.30600000 0.16300000 ;
    END
  END E

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.36900000 0.02700000 0.41400000 0.04500000 ;
        RECT 0.39600000 0.04500000 0.41400000 0.18900000 ;
        RECT 0.36900000 0.18900000 0.41400000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.06300000 0.36000000 0.08100000 ;
      RECT 0.34200000 0.08100000 0.36000000 0.14400000 ;
      RECT 0.01800000 0.08100000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
  END

END OR5x1_ASAP7_75t_L
MACRO XNOR2x2_ASAP7_75t_L
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XNOR2X2_ASAP7_75T_L 0 0 ;
 SIZE  0.5940000000000002 BY 0.2700000000000001 ;
 SYMMETRY X Y ;
 SITE asap7sc7p5t ;
  PIN VSS
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 -0.00900000 0.59400000 0.00900000 ;
    END
  END VSS

  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
       LAYER M1 ;
        RECT 0.00000000 0.26100000 0.59400000 0.27900000 ;
    END
  END VDD

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.12600000 0.12600000 0.14400000 0.18900000 ;
        RECT 0.12600000 0.18900000 0.25200000 0.20700000 ;
        RECT 0.39600000 0.12600000 0.41400000 0.18900000 ;
        RECT 0.34200000 0.18900000 0.41400000 0.20700000 ;
       LAYER M2 ;
        RECT 0.23200000 0.18900000 0.36200000 0.20700000 ;
       LAYER V1 ;
        RECT 0.23200000 0.18900000 0.25000000 0.20700000 ;
        RECT 0.34400000 0.18900000 0.36200000 0.20700000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.18000000 0.12600000 0.19800000 0.14400000 ;
        RECT 0.18000000 0.14400000 0.25200000 0.16200000 ;
        RECT 0.34200000 0.12600000 0.36000000 0.16400000 ;
       LAYER M2 ;
        RECT 0.23200000 0.14400000 0.36000000 0.16200000 ;
       LAYER V1 ;
        RECT 0.23200000 0.14400000 0.25000000 0.16200000 ;
        RECT 0.34200000 0.14400000 0.36000000 0.16200000 ;
    END
  END B

  PIN Y
   DIRECTION OUTPUT ;
   USE SIGNAL ;
    PORT
       LAYER M1 ;
        RECT 0.47700000 0.02700000 0.52200000 0.04500000 ;
        RECT 0.50400000 0.04500000 0.52200000 0.18900000 ;
        RECT 0.47700000 0.18900000 0.52200000 0.20700000 ;
    END
  END Y

  OBS
     LAYER M1 ;
      RECT 0.01800000 0.02700000 0.44100000 0.04500000 ;
      RECT 0.42300000 0.04500000 0.44100000 0.06300000 ;
      RECT 0.42300000 0.06300000 0.46800000 0.08100000 ;
      RECT 0.45000000 0.08100000 0.46800000 0.14400000 ;
      RECT 0.01800000 0.04500000 0.03600000 0.18900000 ;
      RECT 0.01800000 0.18900000 0.06300000 0.20700000 ;
      RECT 0.09900000 0.22500000 0.22500000 0.24300000 ;
      RECT 0.07200000 0.06300000 0.38700000 0.08100000 ;
      RECT 0.07200000 0.08100000 0.09000000 0.14400000 ;
      RECT 0.28800000 0.08100000 0.30600000 0.22500000 ;
      RECT 0.28800000 0.22500000 0.33300000 0.24300000 ;
  END

END XNOR2x2_ASAP7_75t_L
